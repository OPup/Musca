
//------> ./rtl_mgc_ioport.v 
//------------------------------------------------------------------
//                M G C _ I O P O R T _ C O M P S
//------------------------------------------------------------------

//------------------------------------------------------------------
//                       M O D U L E S
//------------------------------------------------------------------

//------------------------------------------------------------------
//-- INPUT ENTITIES
//------------------------------------------------------------------

module mgc_in_wire (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output [width-1:0] d;
  output             lz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule
//------------------------------------------------------------------

module mgc_chan_in (ld, vd, d, lz, vz, z, size, req_size, sizez, sizelz);

  parameter integer rscid = 1;
  parameter integer width = 8;
  parameter integer sz_width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;
  output [sz_width-1:0] size;
  input              req_size;
  input  [sz_width-1:0] sizez;
  output             sizelz;


  wire               vd;
  wire   [width-1:0] d;
  wire               lz;
  wire   [sz_width-1:0] size;
  wire               sizelz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;
  assign size = sizez;
  assign sizelz = req_size;

endmodule


//------------------------------------------------------------------
//-- OUTPUT ENTITIES
//------------------------------------------------------------------

module mgc_out_stdreg (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  input  [width-1:0] d;
  output             lz;
  output [width-1:0] z;

  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_out_prereg_en (ld, d, lz, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    wire               lz;
    wire   [width-1:0] z;

    assign z = d;
    assign lz = ld;

endmodule

//------------------------------------------------------------------
//-- INOUT ENTITIES
//------------------------------------------------------------------

module mgc_inout_stdreg_en (ldin, din, ldout, dout, lzin, lzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    output             lzin;
    output             lzout;
    inout  [width-1:0] z;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign z = ldout ? dout : {width{1'bz}};

endmodule

//------------------------------------------------------------------
module hid_tribuf( I_SIG, ENABLE, O_SIG);
  parameter integer width = 8;

  input [width-1:0] I_SIG;
  input ENABLE;
  inout [width-1:0] O_SIG;

  assign O_SIG = (ENABLE) ? I_SIG : { width{1'bz}};

endmodule
//------------------------------------------------------------------

module mgc_inout_stdreg_wait (ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;
    wire   ldout_and_vzout;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign vdout = vzout ;
    assign ldout_and_vzout = ldout && vzout ;

    hid_tribuf #(width) tb( .I_SIG(dout),
                            .ENABLE(ldout_and_vzout),
                            .O_SIG(z) );

endmodule

//------------------------------------------------------------------

module mgc_inout_buf_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    hid_tribuf #(width) tb( .I_SIG(z_buf),
                            .ENABLE((lzout_buf && (!ldin) && vzout) ),
                            .O_SIG(z)  );

    mgc_out_buf_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFF
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );


endmodule

module mgc_inout_fifo_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer ph_log2 = 3;     // log2(fifo_sz)
    parameter integer pwropt  = 0;     // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               comb;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    assign comb = (lzout_buf && (!ldin) && vzout);

    hid_tribuf #(width) tb2( .I_SIG(z_buf), .ENABLE(comb), .O_SIG(z)  );

    mgc_out_fifo_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
    )
    FIFO
    (
        .clk   (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );

endmodule

//------------------------------------------------------------------
//-- I/O SYNCHRONIZATION ENTITIES
//------------------------------------------------------------------

module mgc_io_sync (ld, lz);

    input  ld;
    output lz;

    assign lz = ld;

endmodule

module mgc_bsync_rdy (rd, rz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 0;

    input  rd;
    output rz;

    wire   rz;

    assign rz = rd;

endmodule

module mgc_bsync_vld (vd, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 0;
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule

module mgc_bsync_rv (rd, vd, rz, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 1;

    input  rd;
    output vd;
    output rz;
    input  vz;

    wire   vd;
    wire   rz;

    assign rz = rd;
    assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_sync (ldin, vdin, ldout, vdout);

  input  ldin;
  output vdin;
  input  ldout;
  output vdout;

  wire   vdin;
  wire   vdout;

  assign vdin = ldout;
  assign vdout = ldin;

endmodule

///////////////////////////////////////////////////////////////////////////////
// dummy function used to preserve funccalls for modulario
// it looks like a memory read to the caller
///////////////////////////////////////////////////////////////////////////////
module funccall_inout (d, ad, bd, z, az, bz);

  parameter integer ram_id = 1;
  parameter integer width = 8;
  parameter integer addr_width = 8;

  output [width-1:0]       d;
  input  [addr_width-1:0]  ad;
  input                    bd;
  input  [width-1:0]       z;
  output [addr_width-1:0]  az;
  output                   bz;

  wire   [width-1:0]       d;
  wire   [addr_width-1:0]  az;
  wire                     bz;

  assign d  = z;
  assign az = ad;
  assign bz = bd;

endmodule


///////////////////////////////////////////////////////////////////////////////
// inlinable modular io not otherwise found in mgc_ioport
///////////////////////////////////////////////////////////////////////////////

module modulario_en_in (vd, d, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output             vd;
  output [width-1:0] d;
  input              vz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               vd;

  assign d = z;
  assign vd = vz;

endmodule

//------> ./rtl_mgc_ioport_v2001.v 
//------------------------------------------------------------------

module mgc_out_reg_pos (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(posedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(posedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg_neg (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(negedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(negedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg (clk, en, arst, srst, ld, d, lz, z); // Not Supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;


    generate
    if (ph_clk == 1'b0)
    begin: NEG_EDGE

        mgc_out_reg_neg
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_neg_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    else
    begin: POS_EDGE

        mgc_out_reg_pos
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_pos_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    endgenerate

endmodule




//------------------------------------------------------------------

module mgc_out_buf_wait (clk, en, arst, srst, ld, vd, d, vz, lz, z); // Not supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    output             vd;
    input  [width-1:0] d;
    output             lz;
    input              vz;
    output [width-1:0] z;

    wire               filled;
    wire               filled_next;
    wire   [width-1:0] abuf;
    wire               lbuf;


    assign filled_next = (filled & (~vz)) | (filled & ld) | (ld & (~vz));

    assign lbuf = ld & ~(filled ^ vz);

    assign vd = vz | ~filled;

    assign lz = ld | filled;

    assign z = (filled) ? abuf : d;

    wire dummy;
    wire dummy_bufreg_lz;

    // Output registers:
    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (1'b1),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    STATREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (filled_next),
        .d       (1'b0),       // input d is unused
        .lz      (filled),
        .z       (dummy)            // output z is unused
    );

    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (lbuf),
        .d       (d),
        .lz      (dummy_bufreg_lz),
        .z       (abuf)
    );

endmodule

//------------------------------------------------------------------

module mgc_out_fifo_wait (clk, en, arst, srst, ld, vd, d, lz, vz,  z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1; // clock enable polarity
    parameter         ph_arst = 1'b1; // async reset polarity
    parameter         ph_srst = 1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt


    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;

    wire    [31:0]      size;


      // Output registers:
 mgc_out_fifo_wait_core#(
        .rscid   (rscid),
        .width   (width),
        .sz_width (32),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
        ) CORE (
        .clk (clk),
        .en (en),
        .arst (arst),
        .srst (srst),
        .ld (ld),
        .vd (vd),
        .d (d),
        .lz (lz),
        .vz (vz),
        .z (z),
        .size (size)
        );

endmodule



module mgc_out_fifo_wait_core (clk, en, arst, srst, ld, vd, d, lz, vz,  z, size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // size of port for elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt

   localparam integer  fifo_b = width * fifo_sz;

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;
    output    [sz_width-1:0]      size;

    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat_pre;
    wire     [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] en_l;
    reg      [(((fifo_sz > 0) ? fifo_sz : 1)-1)/8:0] en_l_s;

    reg       [width-1:0] buff_nxt;

    reg                   stat_nxt;
    reg                   stat_before;
    reg                   stat_after;
    reg                   en_l_var;

    integer               i;
    genvar                eni;

    wire [32:0]           size_t;
    reg [31:0]            count;
    reg [31:0]            count_t;
    reg [32:0]            n_elem;
// pragma translate_off
    reg [31:0]            peak;
// pragma translate_on

    wire [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] dummy_statreg_lz;
    wire [( (fifo_b > 0) ? fifo_b : 1)-1:0] dummy_bufreg_lz;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      assign vd = vz | ~stat[0];
      assign lz = ld | stat[fifo_sz-1];
      assign size_t = (count - (vz && stat[fifo_sz-1])) + ld;
      assign size = size_t[sz_width-1:0];
      assign z = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : d;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          if (i != 0)
            stat_before = stat[i-1];
          else
            stat_before = 1'b0;

          if (i != (fifo_sz-1))
            stat_after = stat[i+1];
          else
            stat_after = 1'b1;

          stat_nxt = stat_after &
                    (stat_before | (stat[i] & (~vz)) | (stat[i] & ld) | (ld & (~vz)));

          stat_pre[i] = stat_nxt;
          en_l_var = 1'b1;
          if (!stat_nxt)
            begin
              buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end
          else if (vz && stat_before)
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
          else if (ld && !((vz && stat_before) || ((!vz) && stat[i])))
            buff_nxt = d;
          else
            begin
              if (pwropt == 0)
                buff_nxt[0+:width] = buff[width*i+:width];
              else
                buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if ((stat_after == 1'b1) && (stat[i] == 1'b0))
            n_elem = ($unsigned(fifo_sz) - 1) - i;
        end

        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b1;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b0;

        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if ((i%'d2) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]|stat_pre[i-1]);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]|stat_pre[i-1]);
          end
        end

        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = { {(32-ph_log2){1'b0}}, fifo_sz};
        else
          count_t = n_elem[31:0];
        count = count_t;
// pragma translate_off
        if ( peak < count )
          peak = count;
// pragma translate_on
      end

      if (pwropt == 0)
      begin: NOCGFIFO
        // Output registers:
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        STATREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
        );
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_b),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        BUFREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre),
            .lz      (dummy_bufreg_lz[0]),
            .z       (buff)
        );
      end
      else
      begin: CGFIFO
        // Output registers:
        if ( pwropt > 1)
        begin: CGSTATFIFO2
          for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
          begin: pwroptGEN1
            mgc_out_reg
            #(
              .rscid   (rscid),
              .width   (1),
              .ph_clk  (ph_clk),
              .ph_en   (ph_en),
              .ph_arst (ph_arst),
              .ph_srst (ph_srst)
            )
            STATREG
            (
              .clk     (clk),
              .en      (en_l_s[eni/8]),
              .arst    (arst),
              .srst    (srst),
              .ld      (1'b1),
              .d       (stat_pre[eni]),
              .lz      (dummy_statreg_lz[eni]),
              .z       (stat[eni])
            );
          end
        end
        else
        begin: CGSTATFIFO
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          STATREG
          (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
          );
        end
        for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
        begin: pwroptGEN2
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (width),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          BUFREG
          (
            .clk     (clk),
            .en      (en_l[eni]),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre[width*eni+:width]),
            .lz      (dummy_bufreg_lz[eni]),
            .z       (buff[width*eni+:width])
          );
        end
      end
    end
    else
    begin: FEED_THRU
      assign vd = vz;
      assign lz = ld;
      assign z = d;
      assign size = ld && !vz;
    end
    endgenerate

endmodule

//------------------------------------------------------------------
//-- PIPE ENTITIES
//------------------------------------------------------------------
/*
 *
 *             _______________________________________________
 * WRITER    |                                               |          READER
 *           |           MGC_PIPE                            |
 *           |           __________________________          |
 *        --<| vdout  --<| vd ---------------  vz<|-----ldin<|---
 *           |           |      FIFO              |          |
 *        ---|>ldout  ---|>ld ---------------- lz |> ---vdin |>--
 *        ---|>dout -----|>d  ---------------- dz |> ----din |>--
 *           |           |________________________|          |
 *           |_______________________________________________|
 */
// two clock pipe
module mgc_pipe (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, size, req_size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer log2_sz = 3; // log2(fifo_sz)
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer pwropt  = 0; // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output [sz_width-1:0]      size;
    input              req_size;


    mgc_out_fifo_wait_core
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz),
        .pwropt   (pwropt)
    )
    FIFO
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (vdin),
        .vz      (ldin),
        .z       (din),
        .size    (size)
    );

endmodule


//------> C:/PROGRA~1/CALYPT~1/CATAPU~1.126/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
         divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
            rmod = {(width_b){1'b0}} - rmod;
         if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2011a.126 Production Release
//  HLS Date:       Wed Aug  8 00:52:07 PDT 2012
// 
//  Generated by:   oh1015@EEWS104A-005
//  Generated date: Wed Apr 27 15:35:15 2016
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    HSVRGB_core
// ------------------------------------------------------------------


module HSVRGB_core (
  clk, rst, R_IN_rsc_mgc_in_wire_d, G_IN_rsc_mgc_in_wire_d, B_IN_rsc_mgc_in_wire_d,
      H_OUT_rsc_mgc_out_stdreg_d, S_OUT_rsc_mgc_out_stdreg_d, V_OUT_rsc_mgc_out_stdreg_d,
      div_mgc_div_a, div_mgc_div_b, div_mgc_div_z, div_mgc_div_1_a, div_mgc_div_1_b,
      div_mgc_div_1_z, div_mgc_div_2_a, div_mgc_div_2_b, div_mgc_div_2_z, div_mgc_div_3_a,
      div_mgc_div_3_b, div_mgc_div_3_z, div_mgc_div_4_a, div_mgc_div_4_b, div_mgc_div_4_z,
      div_mgc_div_5_a, div_mgc_div_5_b, div_mgc_div_5_z, div_mgc_div_6_a, div_mgc_div_6_b,
      div_mgc_div_6_z, div_mgc_div_7_a, div_mgc_div_7_b, div_mgc_div_7_z, div_mgc_div_8_a,
      div_mgc_div_8_b, div_mgc_div_8_z, div_mgc_div_9_a, div_mgc_div_9_b, div_mgc_div_9_z,
      div_mgc_div_10_a, div_mgc_div_10_b, div_mgc_div_10_z, div_mgc_div_11_a, div_mgc_div_11_b,
      div_mgc_div_11_z, div_mgc_div_12_a, div_mgc_div_12_b, div_mgc_div_12_z, div_mgc_div_13_a,
      div_mgc_div_13_b, div_mgc_div_13_z, div_mgc_div_14_a, div_mgc_div_14_b, div_mgc_div_14_z,
      div_mgc_div_15_a, div_mgc_div_15_b, div_mgc_div_15_z, div_mgc_div_16_a, div_mgc_div_16_b,
      div_mgc_div_16_z, div_mgc_div_17_a, div_mgc_div_17_b, div_mgc_div_17_z, div_mgc_div_18_a,
      div_mgc_div_18_b, div_mgc_div_18_z, div_mgc_div_19_a, div_mgc_div_19_b, div_mgc_div_19_z,
      div_mgc_div_20_a, div_mgc_div_20_b, div_mgc_div_20_z, div_mgc_div_21_a, div_mgc_div_21_b,
      div_mgc_div_21_z, div_mgc_div_22_a, div_mgc_div_22_b, div_mgc_div_22_z, div_mgc_div_23_a,
      div_mgc_div_23_b, div_mgc_div_23_z, div_mgc_div_24_a, div_mgc_div_24_b, div_mgc_div_24_z,
      div_mgc_div_25_a, div_mgc_div_25_b, div_mgc_div_25_z, div_mgc_div_26_a, div_mgc_div_26_b,
      div_mgc_div_26_z, div_mgc_div_27_a, div_mgc_div_27_b, div_mgc_div_27_z, div_mgc_div_28_a,
      div_mgc_div_28_b, div_mgc_div_28_z, div_mgc_div_29_a, div_mgc_div_29_b, div_mgc_div_29_z,
      div_mgc_div_30_a, div_mgc_div_30_b, div_mgc_div_30_z, div_mgc_div_31_a, div_mgc_div_31_b,
      div_mgc_div_31_z, div_mgc_div_32_a, div_mgc_div_32_b, div_mgc_div_32_z, div_mgc_div_33_a,
      div_mgc_div_33_b, div_mgc_div_33_z, div_mgc_div_34_a, div_mgc_div_34_b, div_mgc_div_34_z,
      div_mgc_div_35_a, div_mgc_div_35_b, div_mgc_div_35_z
);
  input clk;
  input rst;
  input [31:0] R_IN_rsc_mgc_in_wire_d;
  input [31:0] G_IN_rsc_mgc_in_wire_d;
  input [31:0] B_IN_rsc_mgc_in_wire_d;
  output [31:0] H_OUT_rsc_mgc_out_stdreg_d;
  reg [31:0] H_OUT_rsc_mgc_out_stdreg_d;
  output [31:0] S_OUT_rsc_mgc_out_stdreg_d;
  reg [31:0] S_OUT_rsc_mgc_out_stdreg_d;
  output [31:0] V_OUT_rsc_mgc_out_stdreg_d;
  reg [31:0] V_OUT_rsc_mgc_out_stdreg_d;
  output [48:0] div_mgc_div_a;
  output [31:0] div_mgc_div_b;
  input [48:0] div_mgc_div_z;
  output [48:0] div_mgc_div_1_a;
  output [31:0] div_mgc_div_1_b;
  input [48:0] div_mgc_div_1_z;
  output [48:0] div_mgc_div_2_a;
  output [31:0] div_mgc_div_2_b;
  input [48:0] div_mgc_div_2_z;
  output [48:0] div_mgc_div_3_a;
  output [31:0] div_mgc_div_3_b;
  input [48:0] div_mgc_div_3_z;
  output [48:0] div_mgc_div_4_a;
  output [31:0] div_mgc_div_4_b;
  input [48:0] div_mgc_div_4_z;
  output [48:0] div_mgc_div_5_a;
  output [31:0] div_mgc_div_5_b;
  input [48:0] div_mgc_div_5_z;
  output [48:0] div_mgc_div_6_a;
  output [31:0] div_mgc_div_6_b;
  input [48:0] div_mgc_div_6_z;
  output [48:0] div_mgc_div_7_a;
  output [31:0] div_mgc_div_7_b;
  input [48:0] div_mgc_div_7_z;
  output [48:0] div_mgc_div_8_a;
  output [31:0] div_mgc_div_8_b;
  input [48:0] div_mgc_div_8_z;
  output [48:0] div_mgc_div_9_a;
  output [31:0] div_mgc_div_9_b;
  input [48:0] div_mgc_div_9_z;
  output [48:0] div_mgc_div_10_a;
  output [31:0] div_mgc_div_10_b;
  input [48:0] div_mgc_div_10_z;
  output [48:0] div_mgc_div_11_a;
  output [31:0] div_mgc_div_11_b;
  input [48:0] div_mgc_div_11_z;
  output [48:0] div_mgc_div_12_a;
  output [31:0] div_mgc_div_12_b;
  input [48:0] div_mgc_div_12_z;
  output [48:0] div_mgc_div_13_a;
  output [31:0] div_mgc_div_13_b;
  input [48:0] div_mgc_div_13_z;
  output [48:0] div_mgc_div_14_a;
  output [31:0] div_mgc_div_14_b;
  input [48:0] div_mgc_div_14_z;
  output [48:0] div_mgc_div_15_a;
  output [31:0] div_mgc_div_15_b;
  input [48:0] div_mgc_div_15_z;
  output [48:0] div_mgc_div_16_a;
  output [31:0] div_mgc_div_16_b;
  input [48:0] div_mgc_div_16_z;
  output [48:0] div_mgc_div_17_a;
  output [31:0] div_mgc_div_17_b;
  input [48:0] div_mgc_div_17_z;
  output [48:0] div_mgc_div_18_a;
  output [31:0] div_mgc_div_18_b;
  input [48:0] div_mgc_div_18_z;
  output [48:0] div_mgc_div_19_a;
  output [31:0] div_mgc_div_19_b;
  input [48:0] div_mgc_div_19_z;
  output [48:0] div_mgc_div_20_a;
  output [31:0] div_mgc_div_20_b;
  input [48:0] div_mgc_div_20_z;
  output [48:0] div_mgc_div_21_a;
  output [31:0] div_mgc_div_21_b;
  input [48:0] div_mgc_div_21_z;
  output [48:0] div_mgc_div_22_a;
  output [31:0] div_mgc_div_22_b;
  input [48:0] div_mgc_div_22_z;
  output [48:0] div_mgc_div_23_a;
  output [31:0] div_mgc_div_23_b;
  input [48:0] div_mgc_div_23_z;
  output [48:0] div_mgc_div_24_a;
  output [31:0] div_mgc_div_24_b;
  input [48:0] div_mgc_div_24_z;
  output [48:0] div_mgc_div_25_a;
  output [31:0] div_mgc_div_25_b;
  input [48:0] div_mgc_div_25_z;
  output [48:0] div_mgc_div_26_a;
  output [31:0] div_mgc_div_26_b;
  input [48:0] div_mgc_div_26_z;
  output [47:0] div_mgc_div_27_a;
  output [31:0] div_mgc_div_27_b;
  input [47:0] div_mgc_div_27_z;
  output [47:0] div_mgc_div_28_a;
  output [31:0] div_mgc_div_28_b;
  input [47:0] div_mgc_div_28_z;
  output [47:0] div_mgc_div_29_a;
  output [31:0] div_mgc_div_29_b;
  input [47:0] div_mgc_div_29_z;
  output [47:0] div_mgc_div_30_a;
  output [31:0] div_mgc_div_30_b;
  input [47:0] div_mgc_div_30_z;
  output [47:0] div_mgc_div_31_a;
  output [31:0] div_mgc_div_31_b;
  input [47:0] div_mgc_div_31_z;
  output [47:0] div_mgc_div_32_a;
  output [31:0] div_mgc_div_32_b;
  input [47:0] div_mgc_div_32_z;
  output [47:0] div_mgc_div_33_a;
  output [31:0] div_mgc_div_33_b;
  input [47:0] div_mgc_div_33_z;
  output [47:0] div_mgc_div_34_a;
  output [31:0] div_mgc_div_34_b;
  input [47:0] div_mgc_div_34_z;
  output [47:0] div_mgc_div_35_a;
  output [31:0] div_mgc_div_35_b;
  input [47:0] div_mgc_div_35_z;


  // Interconnect Declarations
  wire [3:0] else_7_if_1_acc_tmp;
  wire [4:0] nl_else_7_if_1_acc_tmp;
  wire [3:0] else_7_else_1_if_acc_tmp;
  wire [4:0] nl_else_7_else_1_if_acc_tmp;
  wire [3:0] else_7_else_1_else_acc_tmp;
  wire [4:0] nl_else_7_else_1_else_acc_tmp;
  wire else_7_else_1_equal_tmp;
  wire else_7_equal_tmp;
  wire [3:0] else_7_if_acc_tmp;
  wire [4:0] nl_else_7_if_acc_tmp;
  wire if_7_equal_tmp;
  wire [15:0] mux1h_81_tmp;
  wire and_dcpl_15;
  wire and_dcpl_17;
  wire and_dcpl_27;
  wire and_dcpl_124;
  wire and_dcpl_136;
  wire and_dcpl_234;
  wire and_dcpl_235;
  wire and_dcpl_248;
  wire and_dcpl_262;
  wire and_dcpl_276;
  wire and_dcpl_291;
  wire and_dcpl_363;
  wire and_dcpl_364;
  wire and_dcpl_377;
  wire and_dcpl_391;
  wire and_dcpl_405;
  wire and_dcpl_420;
  wire and_dcpl_496;
  wire and_dcpl_508;
  wire and_dcpl_606;
  wire and_dcpl_607;
  wire and_dcpl_620;
  wire and_dcpl_634;
  wire and_dcpl_648;
  wire and_dcpl_663;
  wire and_dcpl_735;
  wire and_dcpl_736;
  wire and_dcpl_749;
  wire and_dcpl_763;
  wire and_dcpl_777;
  wire and_dcpl_792;
  wire and_dcpl_868;
  wire and_dcpl_892;
  wire and_dcpl_916;
  wire and_dcpl_940;
  wire and_dcpl_978;
  wire and_dcpl_979;
  wire and_dcpl_992;
  wire and_dcpl_1006;
  wire and_dcpl_1020;
  wire and_dcpl_1035;
  wire and_dcpl_1107;
  wire and_dcpl_1108;
  wire and_dcpl_1121;
  wire and_dcpl_1135;
  wire and_dcpl_1149;
  wire and_dcpl_1164;
  wire and_dcpl_1240;
  wire and_dcpl_1252;
  wire and_dcpl_1350;
  wire and_dcpl_1351;
  wire and_dcpl_1364;
  wire and_dcpl_1378;
  wire and_dcpl_1392;
  wire and_dcpl_1407;
  wire and_dcpl_1479;
  wire and_dcpl_1480;
  wire and_dcpl_1493;
  wire and_dcpl_1507;
  wire and_dcpl_1521;
  wire and_dcpl_1536;
  wire and_dcpl_1612;
  wire and_dcpl_1636;
  wire and_dcpl_1722;
  wire and_dcpl_1723;
  wire and_dcpl_1737;
  wire and_dcpl_1750;
  wire and_dcpl_1778;
  wire and_dcpl_1806;
  wire and_dcpl_1851;
  wire and_dcpl_1852;
  wire and_dcpl_1865;
  wire and_dcpl_1879;
  wire and_dcpl_1893;
  wire and_dcpl_1908;
  wire and_dcpl_1984;
  wire and_dcpl_2008;
  wire and_dcpl_2094;
  wire and_dcpl_2095;
  wire and_dcpl_2108;
  wire and_dcpl_2123;
  wire and_dcpl_2150;
  wire and_dcpl_2164;
  wire and_dcpl_2223;
  wire and_dcpl_2224;
  wire and_dcpl_2237;
  wire and_dcpl_2251;
  wire and_dcpl_2265;
  wire and_dcpl_2280;
  wire and_dcpl_2356;
  wire and_dcpl_2380;
  wire and_dcpl_2741;
  wire and_dcpl_2742;
  wire and_dcpl_2746;
  wire and_dcpl_2749;
  wire and_dcpl_2757;
  wire and_dcpl_2765;
  wire or_tmp_4;
  wire and_dcpl_2777;
  wire and_dcpl_2778;
  wire and_dcpl_2780;
  wire and_dcpl_2783;
  wire and_dcpl_2789;
  wire and_dcpl_2795;
  wire or_dcpl_555;
  wire and_dcpl_2831;
  wire and_dcpl_2832;
  wire and_dcpl_2835;
  wire and_dcpl_2837;
  wire and_dcpl_2843;
  wire and_dcpl_2849;
  wire and_dcpl_2859;
  wire and_dcpl_2860;
  wire and_dcpl_2863;
  wire and_dcpl_2865;
  wire and_dcpl_2871;
  wire and_dcpl_2877;
  wire and_dcpl_2914;
  wire and_dcpl_2915;
  wire and_dcpl_2916;
  wire and_dcpl_2917;
  wire and_dcpl_2924;
  wire and_dcpl_2934;
  wire and_dcpl_2944;
  wire or_dcpl_564;
  wire and_dcpl_2960;
  wire and_dcpl_2961;
  wire and_dcpl_2963;
  wire and_dcpl_2966;
  wire and_dcpl_2969;
  wire and_dcpl_2973;
  wire and_dcpl_2993;
  wire and_dcpl_3052;
  wire and_dcpl_3053;
  wire and_dcpl_3056;
  wire and_dcpl_3058;
  wire and_dcpl_3064;
  wire and_dcpl_3070;
  wire and_dcpl_3085;
  wire and_dcpl_3144;
  wire and_dcpl_3145;
  wire and_dcpl_3146;
  wire and_dcpl_3149;
  wire and_dcpl_3150;
  wire and_dcpl_3152;
  wire or_tmp_6;
  wire or_tmp_7;
  wire not_tmp_146;
  wire and_dcpl_3155;
  wire and_dcpl_3156;
  wire and_dcpl_3158;
  wire or_tmp_9;
  wire or_tmp_10;
  wire or_tmp_12;
  wire and_tmp;
  wire and_dcpl_3161;
  wire and_dcpl_3162;
  wire and_dcpl_3164;
  wire or_tmp_15;
  wire and_tmp_1;
  wire and_dcpl_3167;
  wire and_dcpl_3168;
  wire and_dcpl_3170;
  wire or_tmp_23;
  wire or_tmp_28;
  wire or_tmp_30;
  wire or_tmp_31;
  wire and_dcpl_3173;
  wire and_dcpl_3174;
  wire and_dcpl_3176;
  wire or_tmp_33;
  wire or_tmp_34;
  wire and_dcpl_3179;
  wire and_dcpl_3180;
  wire and_dcpl_3182;
  wire or_tmp_45;
  wire or_tmp_46;
  wire or_tmp_47;
  wire or_tmp_58;
  wire and_dcpl_3186;
  wire and_dcpl_3188;
  wire or_tmp_60;
  wire or_tmp_64;
  wire or_tmp_74;
  wire and_tmp_14;
  wire or_tmp_79;
  wire and_tmp_22;
  wire mux_tmp_20;
  wire or_tmp_92;
  wire or_tmp_94;
  wire and_dcpl_3238;
  wire and_dcpl_3249;
  wire or_tmp_184;
  wire and_tmp_46;
  wire and_dcpl_3258;
  wire and_tmp_47;
  wire and_dcpl_3264;
  wire or_tmp_206;
  wire and_dcpl_3270;
  wire and_dcpl_3276;
  wire or_tmp_221;
  wire and_dcpl_3280;
  wire and_tmp_60;
  wire and_tmp_68;
  wire mux_tmp_49;
  wire and_dcpl_3332;
  wire and_dcpl_3337;
  wire and_dcpl_3343;
  wire or_tmp_359;
  wire and_tmp_92;
  wire and_dcpl_3350;
  wire and_tmp_93;
  wire and_dcpl_3356;
  wire or_tmp_381;
  wire and_dcpl_3362;
  wire and_dcpl_3368;
  wire or_tmp_396;
  wire and_dcpl_3374;
  wire and_tmp_106;
  wire and_tmp_114;
  wire mux_tmp_78;
  wire and_dcpl_3426;
  wire and_dcpl_3437;
  wire or_tmp_534;
  wire and_tmp_138;
  wire and_tmp_139;
  wire or_tmp_556;
  wire or_tmp_571;
  wire and_dcpl_3468;
  wire and_tmp_152;
  wire and_tmp_160;
  wire mux_tmp_107;
  wire and_dcpl_3522;
  wire and_dcpl_3525;
  wire or_tmp_709;
  wire and_tmp_184;
  wire and_dcpl_3538;
  wire and_tmp_185;
  wire and_dcpl_3544;
  wire or_tmp_731;
  wire and_dcpl_3550;
  wire and_dcpl_3556;
  wire or_tmp_746;
  wire and_dcpl_3564;
  wire and_tmp_198;
  wire and_tmp_206;
  wire mux_tmp_138;
  wire or_tmp_884;
  wire and_tmp_230;
  wire and_tmp_231;
  wire or_tmp_906;
  wire or_tmp_921;
  wire and_tmp_244;
  wire and_tmp_252;
  wire mux_tmp_167;
  wire and_dcpl_3713;
  wire or_tmp_1059;
  wire and_tmp_276;
  wire and_dcpl_3726;
  wire and_tmp_277;
  wire and_dcpl_3732;
  wire or_tmp_1081;
  wire and_dcpl_3738;
  wire and_dcpl_3744;
  wire or_tmp_1096;
  wire and_tmp_290;
  wire and_tmp_298;
  wire mux_tmp_196;
  wire or_tmp_1234;
  wire and_tmp_322;
  wire and_tmp_323;
  wire or_tmp_1256;
  wire or_tmp_1271;
  wire and_tmp_344;
  wire mux_tmp_225;
  wire or_tmp_1409;
  wire mux_tmp_246;
  wire or_tmp_1422;
  wire mux_tmp_248;
  wire or_tmp_1434;
  wire or_tmp_1449;
  wire and_tmp_380;
  wire and_tmp_388;
  wire mux_tmp_258;
  wire and_dcpl_3990;
  wire and_dcpl_3991;
  wire and_dcpl_3992;
  wire and_dcpl_3993;
  wire and_dcpl_3996;
  wire and_dcpl_3997;
  wire and_dcpl_3998;
  wire or_dcpl_854;
  wire or_dcpl_855;
  wire or_dcpl_856;
  wire or_dcpl_857;
  wire and_dcpl_4003;
  wire and_dcpl_4006;
  wire and_dcpl_4010;
  wire and_dcpl_4013;
  wire or_tmp_1591;
  wire or_tmp_1592;
  wire or_tmp_1593;
  wire and_dcpl_4017;
  wire and_dcpl_4020;
  wire or_tmp_1595;
  wire and_dcpl_4024;
  wire and_dcpl_4027;
  wire or_tmp_1600;
  wire and_dcpl_4031;
  wire and_dcpl_4034;
  wire or_tmp_1606;
  wire and_dcpl_4038;
  wire and_dcpl_4041;
  wire or_tmp_1613;
  wire and_tmp_421;
  wire and_dcpl_4098;
  wire and_dcpl_4099;
  wire and_dcpl_4104;
  wire or_dcpl_864;
  wire or_dcpl_865;
  wire and_dcpl_4111;
  wire and_dcpl_4121;
  wire or_tmp_1671;
  wire or_tmp_1672;
  wire or_tmp_1673;
  wire and_dcpl_4125;
  wire or_tmp_1675;
  wire or_tmp_1680;
  wire and_dcpl_4139;
  wire or_tmp_1686;
  wire and_dcpl_4146;
  wire or_tmp_1693;
  wire and_tmp_464;
  wire and_dcpl_4209;
  wire and_dcpl_4212;
  wire or_dcpl_877;
  wire and_dcpl_4219;
  wire and_dcpl_4226;
  wire or_tmp_1751;
  wire or_tmp_1752;
  wire or_tmp_1753;
  wire and_dcpl_4233;
  wire or_tmp_1755;
  wire or_tmp_1760;
  wire and_dcpl_4247;
  wire or_tmp_1766;
  wire and_dcpl_4254;
  wire or_tmp_1773;
  wire and_tmp_507;
  wire and_dcpl_4320;
  wire and_dcpl_4327;
  wire or_tmp_1831;
  wire or_tmp_1832;
  wire or_tmp_1833;
  wire and_dcpl_4341;
  wire or_tmp_1835;
  wire or_tmp_1840;
  wire and_dcpl_4355;
  wire or_tmp_1846;
  wire and_dcpl_4362;
  wire or_tmp_1853;
  wire and_tmp_550;
  wire and_dcpl_4423;
  wire and_dcpl_4430;
  wire or_dcpl_895;
  wire and_dcpl_4438;
  wire and_dcpl_4442;
  wire or_tmp_1911;
  wire or_tmp_1912;
  wire or_tmp_1913;
  wire and_dcpl_4452;
  wire or_tmp_1915;
  wire or_tmp_1920;
  wire and_dcpl_4466;
  wire or_tmp_1926;
  wire and_dcpl_4473;
  wire or_tmp_1933;
  wire and_tmp_593;
  wire and_dcpl_4531;
  wire or_dcpl_905;
  wire or_tmp_1991;
  wire or_tmp_1992;
  wire or_tmp_1993;
  wire or_tmp_1995;
  wire or_tmp_2000;
  wire or_tmp_2006;
  wire or_tmp_2013;
  wire and_tmp_636;
  wire and_dcpl_4658;
  wire or_tmp_2071;
  wire or_tmp_2072;
  wire or_tmp_2073;
  wire or_tmp_2075;
  wire or_tmp_2080;
  wire or_tmp_2086;
  wire or_tmp_2093;
  wire and_tmp_679;
  wire or_tmp_2151;
  wire or_tmp_2152;
  wire or_tmp_2153;
  wire or_tmp_2155;
  wire or_tmp_2160;
  wire or_tmp_2166;
  wire or_tmp_2173;
  wire and_tmp_722;
  wire or_dcpl_935;
  wire or_tmp_2231;
  wire or_tmp_2232;
  wire or_tmp_2233;
  wire mux_tmp_376;
  wire or_tmp_2236;
  wire or_tmp_2243;
  wire or_tmp_2252;
  wire and_tmp_755;
  wire mux_tmp_390;
  wire mux_tmp_391;
  wire mux_tmp_392;
  wire and_dcpl_4962;
  wire and_dcpl_4963;
  wire and_dcpl_4965;
  wire and_dcpl_4966;
  wire and_dcpl_4968;
  wire and_dcpl_4969;
  wire and_dcpl_4971;
  wire and_dcpl_4972;
  wire or_dcpl_944;
  wire or_dcpl_945;
  wire or_dcpl_947;
  wire or_dcpl_948;
  wire and_dcpl_4981;
  wire and_dcpl_4989;
  wire or_tmp_2353;
  wire or_tmp_2354;
  wire or_tmp_2355;
  wire and_tmp_760;
  wire and_dcpl_4997;
  wire or_tmp_2360;
  wire and_tmp_762;
  wire and_dcpl_5005;
  wire or_tmp_2363;
  wire and_tmp_763;
  wire and_tmp_765;
  wire and_dcpl_5013;
  wire or_tmp_2369;
  wire and_tmp_769;
  wire and_dcpl_5021;
  wire or_tmp_2376;
  wire and_tmp_774;
  wire and_tmp_780;
  wire and_dcpl_5086;
  wire and_dcpl_5087;
  wire or_dcpl_956;
  wire or_dcpl_957;
  wire or_tmp_2433;
  wire or_tmp_2434;
  wire or_tmp_2435;
  wire and_tmp_803;
  wire or_tmp_2440;
  wire and_tmp_805;
  wire or_tmp_2443;
  wire and_tmp_806;
  wire and_tmp_808;
  wire or_tmp_2449;
  wire and_tmp_812;
  wire or_tmp_2456;
  wire and_tmp_817;
  wire and_tmp_823;
  wire and_dcpl_5214;
  wire and_dcpl_5216;
  wire or_dcpl_972;
  wire or_tmp_2513;
  wire or_tmp_2514;
  wire or_tmp_2515;
  wire and_tmp_846;
  wire or_tmp_2520;
  wire and_tmp_848;
  wire or_tmp_2523;
  wire and_tmp_849;
  wire and_tmp_851;
  wire or_tmp_2529;
  wire and_tmp_855;
  wire or_tmp_2536;
  wire and_tmp_860;
  wire and_tmp_866;
  wire or_tmp_2593;
  wire or_tmp_2594;
  wire or_tmp_2595;
  wire and_tmp_889;
  wire or_tmp_2600;
  wire and_tmp_891;
  wire or_tmp_2603;
  wire and_tmp_892;
  wire and_tmp_894;
  wire or_tmp_2609;
  wire and_tmp_898;
  wire or_tmp_2616;
  wire and_tmp_903;
  wire and_tmp_909;
  wire and_dcpl_5459;
  wire and_dcpl_5464;
  wire or_dcpl_993;
  wire or_tmp_2673;
  wire or_tmp_2674;
  wire or_tmp_2675;
  wire and_tmp_932;
  wire or_tmp_2680;
  wire and_tmp_934;
  wire or_tmp_2683;
  wire and_tmp_935;
  wire and_tmp_937;
  wire or_tmp_2689;
  wire and_tmp_941;
  wire or_tmp_2696;
  wire and_tmp_946;
  wire and_tmp_952;
  wire and_dcpl_5583;
  wire or_dcpl_1005;
  wire or_tmp_2753;
  wire or_tmp_2754;
  wire or_tmp_2755;
  wire and_tmp_975;
  wire or_tmp_2760;
  wire and_tmp_977;
  wire or_tmp_2763;
  wire and_tmp_978;
  wire and_tmp_980;
  wire or_tmp_2769;
  wire and_tmp_984;
  wire or_tmp_2776;
  wire and_tmp_989;
  wire and_tmp_995;
  wire and_dcpl_5712;
  wire or_tmp_2833;
  wire or_tmp_2834;
  wire or_tmp_2835;
  wire and_tmp_1018;
  wire or_tmp_2840;
  wire and_tmp_1020;
  wire or_tmp_2843;
  wire and_tmp_1021;
  wire and_tmp_1023;
  wire or_tmp_2849;
  wire and_tmp_1027;
  wire or_tmp_2856;
  wire and_tmp_1032;
  wire and_tmp_1038;
  wire or_tmp_2913;
  wire or_tmp_2914;
  wire or_tmp_2915;
  wire and_tmp_1061;
  wire or_tmp_2920;
  wire and_tmp_1063;
  wire or_tmp_2923;
  wire and_tmp_1064;
  wire and_tmp_1066;
  wire or_tmp_2929;
  wire and_tmp_1070;
  wire or_tmp_2936;
  wire and_tmp_1075;
  wire and_tmp_1081;
  wire or_dcpl_1041;
  wire or_tmp_2993;
  wire or_tmp_2994;
  wire or_tmp_2995;
  wire or_tmp_2996;
  wire and_tmp_1104;
  wire or_tmp_3001;
  wire and_tmp_1105;
  wire mux_tmp_523;
  wire or_tmp_3006;
  wire mux_tmp_525;
  wire mux_tmp_526;
  wire or_tmp_3015;
  wire or_tmp_3026;
  wire mux_tmp_540;
  wire mux_tmp_541;
  wire mux_tmp_542;
  wire and_tmp_1106;
  wire and_dcpl_6078;
  wire and_dcpl_6079;
  wire and_dcpl_6082;
  wire and_dcpl_6084;
  wire and_dcpl_6085;
  wire and_dcpl_6088;
  wire or_dcpl_1052;
  wire or_dcpl_1053;
  wire or_dcpl_1056;
  wire or_tmp_3115;
  wire or_tmp_3116;
  wire or_tmp_3117;
  wire or_tmp_3121;
  wire or_tmp_3123;
  wire and_tmp_1116;
  wire or_tmp_3128;
  wire or_tmp_3134;
  wire and_dcpl_6202;
  wire and_dcpl_6203;
  wire and_dcpl_6209;
  wire or_dcpl_1064;
  wire or_dcpl_1065;
  wire or_tmp_3183;
  wire or_tmp_3184;
  wire or_tmp_3185;
  wire or_tmp_3189;
  wire or_tmp_3191;
  wire and_tmp_1171;
  wire or_tmp_3196;
  wire or_tmp_3202;
  wire and_dcpl_6330;
  wire and_dcpl_6332;
  wire and_dcpl_6333;
  wire or_dcpl_1080;
  wire or_tmp_3251;
  wire or_tmp_3252;
  wire or_tmp_3253;
  wire or_tmp_3257;
  wire or_tmp_3259;
  wire and_tmp_1226;
  wire or_tmp_3264;
  wire or_tmp_3270;
  wire and_dcpl_6457;
  wire or_tmp_3319;
  wire or_tmp_3320;
  wire or_tmp_3321;
  wire or_tmp_3325;
  wire or_tmp_3327;
  wire and_tmp_1281;
  wire or_tmp_3332;
  wire or_tmp_3338;
  wire and_dcpl_6575;
  wire and_dcpl_6584;
  wire or_dcpl_1101;
  wire or_tmp_3387;
  wire or_tmp_3388;
  wire or_tmp_3389;
  wire or_tmp_3393;
  wire or_tmp_3395;
  wire and_tmp_1336;
  wire or_tmp_3400;
  wire or_tmp_3406;
  wire and_dcpl_6699;
  wire or_dcpl_1113;
  wire or_tmp_3455;
  wire or_tmp_3456;
  wire or_tmp_3457;
  wire or_tmp_3461;
  wire or_tmp_3463;
  wire and_tmp_1391;
  wire or_tmp_3468;
  wire or_tmp_3474;
  wire or_tmp_3523;
  wire or_tmp_3524;
  wire or_tmp_3525;
  wire or_tmp_3529;
  wire or_tmp_3531;
  wire and_tmp_1446;
  wire or_tmp_3536;
  wire or_tmp_3542;
  wire or_tmp_3591;
  wire or_tmp_3592;
  wire or_tmp_3593;
  wire or_tmp_3597;
  wire or_tmp_3599;
  wire and_tmp_1501;
  wire or_tmp_3604;
  wire or_tmp_3610;
  wire or_dcpl_1149;
  wire or_tmp_3659;
  wire or_tmp_3660;
  wire or_tmp_3661;
  wire or_tmp_3662;
  wire or_tmp_3666;
  wire and_tmp_1553;
  wire or_tmp_3670;
  wire mux_tmp_571;
  wire mux_tmp_572;
  wire or_tmp_3678;
  wire or_tmp_3688;
  wire mux_tmp_583;
  wire mux_tmp_584;
  wire mux_tmp_585;
  wire or_dcpl_1160;
  wire or_dcpl_1161;
  wire or_dcpl_1162;
  wire or_dcpl_1170;
  wire or_dcpl_1180;
  wire or_dcpl_1190;
  wire or_dcpl_1202;
  reg [15:0] else_7_acc_2_psp_sg1_sva;
  reg [3:0] else_7_if_div_9cyc;
  reg [3:0] else_7_if_1_div_9cyc;
  reg [29:0] h_2_sva_duc;
  reg [3:0] else_7_else_1_if_div_9cyc;
  reg [29:0] div_sdt_2_sva_duc;
  reg [3:0] else_7_else_1_else_div_9cyc;
  reg [29:0] div_sdt_3_sva_duc;
  reg else_7_else_1_equal_svs_1;
  reg if_7_equal_svs_9;
  reg unequal_tmp_1;
  reg unequal_tmp_2;
  reg unequal_tmp_3;
  reg unequal_tmp_4;
  reg unequal_tmp_5;
  reg unequal_tmp_6;
  reg unequal_tmp_7;
  reg unequal_tmp_8;
  reg unequal_tmp_9;
  reg else_7_equal_svs_9;
  reg [3:0] else_7_if_div_9cyc_st;
  reg else_7_and_5_itm_1;
  reg else_7_and_5_itm_2;
  reg else_7_and_5_itm_3;
  reg else_7_and_5_itm_4;
  reg else_7_and_5_itm_5;
  reg else_7_and_5_itm_6;
  reg else_7_and_5_itm_7;
  reg else_7_and_5_itm_8;
  reg else_7_and_5_itm_9;
  reg [14:0] slc_3_itm_1;
  reg [14:0] slc_3_itm_2;
  reg [14:0] slc_3_itm_3;
  reg [14:0] slc_3_itm_4;
  reg [14:0] slc_3_itm_5;
  reg [14:0] slc_3_itm_6;
  reg [14:0] slc_3_itm_7;
  reg [14:0] slc_3_itm_8;
  reg [14:0] slc_3_itm_9;
  reg if_7_equal_svs_st_1;
  reg if_7_equal_svs_st_2;
  reg if_7_equal_svs_st_3;
  reg if_7_equal_svs_st_4;
  reg if_7_equal_svs_st_5;
  reg if_7_equal_svs_st_6;
  reg if_7_equal_svs_st_7;
  reg if_7_equal_svs_st_8;
  reg [15:0] max_sg1_lpi_dfm_3_st_1;
  reg [15:0] max_sg1_lpi_dfm_3_st_2;
  reg [15:0] max_sg1_lpi_dfm_3_st_3;
  reg [15:0] max_sg1_lpi_dfm_3_st_4;
  reg [15:0] max_sg1_lpi_dfm_3_st_5;
  reg [15:0] max_sg1_lpi_dfm_3_st_6;
  reg [15:0] max_sg1_lpi_dfm_3_st_7;
  reg [15:0] max_sg1_lpi_dfm_3_st_8;
  reg [3:0] else_7_if_div_9cyc_st_1;
  reg [3:0] else_7_if_div_9cyc_st_2;
  reg [3:0] else_7_if_div_9cyc_st_3;
  reg [3:0] else_7_if_div_9cyc_st_4;
  reg [3:0] else_7_if_div_9cyc_st_5;
  reg [3:0] else_7_if_div_9cyc_st_6;
  reg [3:0] else_7_if_div_9cyc_st_7;
  reg [3:0] else_7_if_div_9cyc_st_8;
  reg [15:0] max_sg1_lpi_dfm_3_st_9;
  reg [3:0] else_7_if_div_9cyc_st_9;
  reg else_7_equal_svs_st_1;
  reg else_7_equal_svs_st_2;
  reg else_7_equal_svs_st_3;
  reg else_7_equal_svs_st_4;
  reg else_7_equal_svs_st_5;
  reg else_7_equal_svs_st_6;
  reg else_7_equal_svs_st_7;
  reg else_7_equal_svs_st_8;
  reg [3:0] else_7_if_1_div_9cyc_st_2;
  reg [3:0] else_7_if_1_div_9cyc_st_3;
  reg [3:0] else_7_if_1_div_9cyc_st_4;
  reg [3:0] else_7_if_1_div_9cyc_st_5;
  reg [3:0] else_7_if_1_div_9cyc_st_6;
  reg [3:0] else_7_if_1_div_9cyc_st_7;
  reg [3:0] else_7_if_1_div_9cyc_st_8;
  reg [3:0] else_7_if_1_div_9cyc_st_9;
  reg else_7_else_1_equal_svs_st_2;
  reg else_7_else_1_equal_svs_st_3;
  reg else_7_else_1_equal_svs_st_4;
  reg else_7_else_1_equal_svs_st_5;
  reg else_7_else_1_equal_svs_st_6;
  reg else_7_else_1_equal_svs_st_7;
  reg else_7_else_1_equal_svs_st_8;
  reg [3:0] else_7_else_1_if_div_9cyc_st_2;
  reg [3:0] else_7_else_1_if_div_9cyc_st_3;
  reg [3:0] else_7_else_1_if_div_9cyc_st_4;
  reg [3:0] else_7_else_1_if_div_9cyc_st_5;
  reg [3:0] else_7_else_1_if_div_9cyc_st_6;
  reg [3:0] else_7_else_1_if_div_9cyc_st_7;
  reg [3:0] else_7_else_1_if_div_9cyc_st_8;
  reg else_7_else_1_equal_svs_st_9;
  reg [3:0] else_7_else_1_if_div_9cyc_st_9;
  reg [3:0] else_7_else_1_else_div_9cyc_st_2;
  reg [3:0] else_7_else_1_else_div_9cyc_st_3;
  reg [3:0] else_7_else_1_else_div_9cyc_st_4;
  reg [3:0] else_7_else_1_else_div_9cyc_st_5;
  reg [3:0] else_7_else_1_else_div_9cyc_st_6;
  reg [3:0] else_7_else_1_else_div_9cyc_st_7;
  reg [3:0] else_7_else_1_else_div_9cyc_st_8;
  reg [3:0] else_7_else_1_else_div_9cyc_st_9;
  reg main_stage_0_2;
  reg main_stage_0_3;
  reg main_stage_0_4;
  reg main_stage_0_5;
  reg main_stage_0_6;
  reg main_stage_0_7;
  reg main_stage_0_8;
  reg main_stage_0_9;
  reg main_stage_0_10;
  reg [15:0] else_7_if_div_tmp_duc_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_9_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_10_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_11_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_12_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_13_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_14_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_15_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_16_sg1;
  reg [15:0] delta_conc_1_tmp_mut_9_sg1;
  reg [15:0] delta_conc_1_tmp_mut_10_sg1;
  reg [15:0] delta_conc_1_tmp_mut_11_sg1;
  reg [15:0] delta_conc_1_tmp_mut_12_sg1;
  reg [15:0] delta_conc_1_tmp_mut_13_sg1;
  reg [15:0] delta_conc_1_tmp_mut_14_sg1;
  reg [15:0] delta_conc_1_tmp_mut_15_sg1;
  reg [15:0] delta_conc_1_tmp_mut_16_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_9_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_10_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_11_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_12_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_13_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_14_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_15_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_16_sg1;
  reg [15:0] delta_conc_3_tmp_mut_9_sg1;
  reg [15:0] delta_conc_3_tmp_mut_10_sg1;
  reg [15:0] delta_conc_3_tmp_mut_11_sg1;
  reg [15:0] delta_conc_3_tmp_mut_12_sg1;
  reg [15:0] delta_conc_3_tmp_mut_13_sg1;
  reg [15:0] delta_conc_3_tmp_mut_14_sg1;
  reg [15:0] delta_conc_3_tmp_mut_15_sg1;
  reg [15:0] delta_conc_3_tmp_mut_16_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_17_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_18_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_19_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_20_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_21_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_22_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_23_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_24_sg1;
  reg [15:0] delta_conc_3_tmp_mut_17_sg1;
  reg [15:0] delta_conc_3_tmp_mut_18_sg1;
  reg [15:0] delta_conc_3_tmp_mut_19_sg1;
  reg [15:0] delta_conc_3_tmp_mut_20_sg1;
  reg [15:0] delta_conc_3_tmp_mut_21_sg1;
  reg [15:0] delta_conc_3_tmp_mut_22_sg1;
  reg [15:0] delta_conc_3_tmp_mut_23_sg1;
  reg [15:0] delta_conc_3_tmp_mut_24_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_25_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_26_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_27_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_28_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_29_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_30_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_31_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_32_sg1;
  reg [15:0] delta_conc_3_tmp_mut_25_sg1;
  reg [15:0] delta_conc_3_tmp_mut_26_sg1;
  reg [15:0] delta_conc_3_tmp_mut_27_sg1;
  reg [15:0] delta_conc_3_tmp_mut_28_sg1;
  reg [15:0] delta_conc_3_tmp_mut_29_sg1;
  reg [15:0] delta_conc_3_tmp_mut_30_sg1;
  reg [15:0] delta_conc_3_tmp_mut_31_sg1;
  reg [15:0] delta_conc_3_tmp_mut_32_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_33_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_34_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_35_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_36_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_37_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_38_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_39_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_40_sg1;
  reg [15:0] delta_conc_3_tmp_mut_33_sg1;
  reg [15:0] delta_conc_3_tmp_mut_34_sg1;
  reg [15:0] delta_conc_3_tmp_mut_35_sg1;
  reg [15:0] delta_conc_3_tmp_mut_36_sg1;
  reg [15:0] delta_conc_3_tmp_mut_37_sg1;
  reg [15:0] delta_conc_3_tmp_mut_38_sg1;
  reg [15:0] delta_conc_3_tmp_mut_39_sg1;
  reg [15:0] delta_conc_3_tmp_mut_40_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_41_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_42_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_43_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_44_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_45_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_46_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_47_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_48_sg1;
  reg [15:0] delta_conc_3_tmp_mut_41_sg1;
  reg [15:0] delta_conc_3_tmp_mut_42_sg1;
  reg [15:0] delta_conc_3_tmp_mut_43_sg1;
  reg [15:0] delta_conc_3_tmp_mut_44_sg1;
  reg [15:0] delta_conc_3_tmp_mut_45_sg1;
  reg [15:0] delta_conc_3_tmp_mut_46_sg1;
  reg [15:0] delta_conc_3_tmp_mut_47_sg1;
  reg [15:0] delta_conc_3_tmp_mut_48_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_49_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_50_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_51_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_52_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_53_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_54_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_55_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_56_sg1;
  reg [15:0] delta_conc_3_tmp_mut_49_sg1;
  reg [15:0] delta_conc_3_tmp_mut_50_sg1;
  reg [15:0] delta_conc_3_tmp_mut_51_sg1;
  reg [15:0] delta_conc_3_tmp_mut_52_sg1;
  reg [15:0] delta_conc_3_tmp_mut_53_sg1;
  reg [15:0] delta_conc_3_tmp_mut_54_sg1;
  reg [15:0] delta_conc_3_tmp_mut_55_sg1;
  reg [15:0] delta_conc_3_tmp_mut_56_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_57_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_58_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_59_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_60_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_61_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_62_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_63_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_64_sg1;
  reg [15:0] delta_conc_3_tmp_mut_57_sg1;
  reg [15:0] delta_conc_3_tmp_mut_58_sg1;
  reg [15:0] delta_conc_3_tmp_mut_59_sg1;
  reg [15:0] delta_conc_3_tmp_mut_60_sg1;
  reg [15:0] delta_conc_3_tmp_mut_61_sg1;
  reg [15:0] delta_conc_3_tmp_mut_62_sg1;
  reg [15:0] delta_conc_3_tmp_mut_63_sg1;
  reg [15:0] delta_conc_3_tmp_mut_64_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_65_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_66_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_67_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_68_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_69_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_70_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_71_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_72_sg1;
  reg [15:0] delta_conc_3_tmp_mut_65_sg1;
  reg [15:0] delta_conc_3_tmp_mut_66_sg1;
  reg [15:0] delta_conc_3_tmp_mut_67_sg1;
  reg [15:0] delta_conc_3_tmp_mut_68_sg1;
  reg [15:0] delta_conc_3_tmp_mut_69_sg1;
  reg [15:0] delta_conc_3_tmp_mut_70_sg1;
  reg [15:0] delta_conc_3_tmp_mut_71_sg1;
  reg [15:0] delta_conc_3_tmp_mut_72_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_73_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_74_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_75_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_76_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_77_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_78_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_79_sg1;
  reg [16:0] else_7_else_1_else_conc_tmp_mut_80_sg1;
  reg [15:0] delta_conc_3_tmp_mut_73_sg1;
  reg [15:0] delta_conc_3_tmp_mut_74_sg1;
  reg [15:0] delta_conc_3_tmp_mut_75_sg1;
  reg [15:0] delta_conc_3_tmp_mut_76_sg1;
  reg [15:0] delta_conc_3_tmp_mut_77_sg1;
  reg [15:0] delta_conc_3_tmp_mut_78_sg1;
  reg [15:0] delta_conc_3_tmp_mut_79_sg1;
  reg [15:0] delta_conc_3_tmp_mut_80_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_9_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_10_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_11_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_12_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_13_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_14_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_15_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_16_sg1;
  reg [15:0] delta_conc_2_tmp_mut_9_sg1;
  reg [15:0] delta_conc_2_tmp_mut_10_sg1;
  reg [15:0] delta_conc_2_tmp_mut_11_sg1;
  reg [15:0] delta_conc_2_tmp_mut_12_sg1;
  reg [15:0] delta_conc_2_tmp_mut_13_sg1;
  reg [15:0] delta_conc_2_tmp_mut_14_sg1;
  reg [15:0] delta_conc_2_tmp_mut_15_sg1;
  reg [15:0] delta_conc_2_tmp_mut_16_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_17_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_18_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_19_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_20_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_21_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_22_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_23_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_24_sg1;
  reg [15:0] delta_conc_2_tmp_mut_17_sg1;
  reg [15:0] delta_conc_2_tmp_mut_18_sg1;
  reg [15:0] delta_conc_2_tmp_mut_19_sg1;
  reg [15:0] delta_conc_2_tmp_mut_20_sg1;
  reg [15:0] delta_conc_2_tmp_mut_21_sg1;
  reg [15:0] delta_conc_2_tmp_mut_22_sg1;
  reg [15:0] delta_conc_2_tmp_mut_23_sg1;
  reg [15:0] delta_conc_2_tmp_mut_24_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_25_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_26_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_27_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_28_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_29_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_30_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_31_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_32_sg1;
  reg [15:0] delta_conc_2_tmp_mut_25_sg1;
  reg [15:0] delta_conc_2_tmp_mut_26_sg1;
  reg [15:0] delta_conc_2_tmp_mut_27_sg1;
  reg [15:0] delta_conc_2_tmp_mut_28_sg1;
  reg [15:0] delta_conc_2_tmp_mut_29_sg1;
  reg [15:0] delta_conc_2_tmp_mut_30_sg1;
  reg [15:0] delta_conc_2_tmp_mut_31_sg1;
  reg [15:0] delta_conc_2_tmp_mut_32_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_33_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_34_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_35_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_36_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_37_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_38_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_39_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_40_sg1;
  reg [15:0] delta_conc_2_tmp_mut_33_sg1;
  reg [15:0] delta_conc_2_tmp_mut_34_sg1;
  reg [15:0] delta_conc_2_tmp_mut_35_sg1;
  reg [15:0] delta_conc_2_tmp_mut_36_sg1;
  reg [15:0] delta_conc_2_tmp_mut_37_sg1;
  reg [15:0] delta_conc_2_tmp_mut_38_sg1;
  reg [15:0] delta_conc_2_tmp_mut_39_sg1;
  reg [15:0] delta_conc_2_tmp_mut_40_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_41_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_42_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_43_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_44_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_45_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_46_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_47_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_48_sg1;
  reg [15:0] delta_conc_2_tmp_mut_41_sg1;
  reg [15:0] delta_conc_2_tmp_mut_42_sg1;
  reg [15:0] delta_conc_2_tmp_mut_43_sg1;
  reg [15:0] delta_conc_2_tmp_mut_44_sg1;
  reg [15:0] delta_conc_2_tmp_mut_45_sg1;
  reg [15:0] delta_conc_2_tmp_mut_46_sg1;
  reg [15:0] delta_conc_2_tmp_mut_47_sg1;
  reg [15:0] delta_conc_2_tmp_mut_48_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_49_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_50_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_51_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_52_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_53_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_54_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_55_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_56_sg1;
  reg [15:0] delta_conc_2_tmp_mut_49_sg1;
  reg [15:0] delta_conc_2_tmp_mut_50_sg1;
  reg [15:0] delta_conc_2_tmp_mut_51_sg1;
  reg [15:0] delta_conc_2_tmp_mut_52_sg1;
  reg [15:0] delta_conc_2_tmp_mut_53_sg1;
  reg [15:0] delta_conc_2_tmp_mut_54_sg1;
  reg [15:0] delta_conc_2_tmp_mut_55_sg1;
  reg [15:0] delta_conc_2_tmp_mut_56_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_57_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_58_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_59_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_60_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_61_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_62_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_63_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_64_sg1;
  reg [15:0] delta_conc_2_tmp_mut_57_sg1;
  reg [15:0] delta_conc_2_tmp_mut_58_sg1;
  reg [15:0] delta_conc_2_tmp_mut_59_sg1;
  reg [15:0] delta_conc_2_tmp_mut_60_sg1;
  reg [15:0] delta_conc_2_tmp_mut_61_sg1;
  reg [15:0] delta_conc_2_tmp_mut_62_sg1;
  reg [15:0] delta_conc_2_tmp_mut_63_sg1;
  reg [15:0] delta_conc_2_tmp_mut_64_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_65_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_66_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_67_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_68_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_69_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_70_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_71_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_72_sg1;
  reg [15:0] delta_conc_2_tmp_mut_65_sg1;
  reg [15:0] delta_conc_2_tmp_mut_66_sg1;
  reg [15:0] delta_conc_2_tmp_mut_67_sg1;
  reg [15:0] delta_conc_2_tmp_mut_68_sg1;
  reg [15:0] delta_conc_2_tmp_mut_69_sg1;
  reg [15:0] delta_conc_2_tmp_mut_70_sg1;
  reg [15:0] delta_conc_2_tmp_mut_71_sg1;
  reg [15:0] delta_conc_2_tmp_mut_72_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_73_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_74_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_75_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_76_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_77_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_78_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_79_sg1;
  reg [16:0] else_7_else_1_if_conc_tmp_mut_80_sg1;
  reg [15:0] delta_conc_2_tmp_mut_73_sg1;
  reg [15:0] delta_conc_2_tmp_mut_74_sg1;
  reg [15:0] delta_conc_2_tmp_mut_75_sg1;
  reg [15:0] delta_conc_2_tmp_mut_76_sg1;
  reg [15:0] delta_conc_2_tmp_mut_77_sg1;
  reg [15:0] delta_conc_2_tmp_mut_78_sg1;
  reg [15:0] delta_conc_2_tmp_mut_79_sg1;
  reg [15:0] delta_conc_2_tmp_mut_80_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_17_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_18_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_19_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_20_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_21_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_22_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_23_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_24_sg1;
  reg [15:0] delta_conc_1_tmp_mut_17_sg1;
  reg [15:0] delta_conc_1_tmp_mut_18_sg1;
  reg [15:0] delta_conc_1_tmp_mut_19_sg1;
  reg [15:0] delta_conc_1_tmp_mut_20_sg1;
  reg [15:0] delta_conc_1_tmp_mut_21_sg1;
  reg [15:0] delta_conc_1_tmp_mut_22_sg1;
  reg [15:0] delta_conc_1_tmp_mut_23_sg1;
  reg [15:0] delta_conc_1_tmp_mut_24_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_25_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_26_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_27_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_28_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_29_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_30_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_31_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_32_sg1;
  reg [15:0] delta_conc_1_tmp_mut_25_sg1;
  reg [15:0] delta_conc_1_tmp_mut_26_sg1;
  reg [15:0] delta_conc_1_tmp_mut_27_sg1;
  reg [15:0] delta_conc_1_tmp_mut_28_sg1;
  reg [15:0] delta_conc_1_tmp_mut_29_sg1;
  reg [15:0] delta_conc_1_tmp_mut_30_sg1;
  reg [15:0] delta_conc_1_tmp_mut_31_sg1;
  reg [15:0] delta_conc_1_tmp_mut_32_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_33_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_34_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_35_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_36_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_37_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_38_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_39_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_40_sg1;
  reg [15:0] delta_conc_1_tmp_mut_33_sg1;
  reg [15:0] delta_conc_1_tmp_mut_34_sg1;
  reg [15:0] delta_conc_1_tmp_mut_35_sg1;
  reg [15:0] delta_conc_1_tmp_mut_36_sg1;
  reg [15:0] delta_conc_1_tmp_mut_37_sg1;
  reg [15:0] delta_conc_1_tmp_mut_38_sg1;
  reg [15:0] delta_conc_1_tmp_mut_39_sg1;
  reg [15:0] delta_conc_1_tmp_mut_40_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_41_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_42_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_43_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_44_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_45_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_46_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_47_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_48_sg1;
  reg [15:0] delta_conc_1_tmp_mut_41_sg1;
  reg [15:0] delta_conc_1_tmp_mut_42_sg1;
  reg [15:0] delta_conc_1_tmp_mut_43_sg1;
  reg [15:0] delta_conc_1_tmp_mut_44_sg1;
  reg [15:0] delta_conc_1_tmp_mut_45_sg1;
  reg [15:0] delta_conc_1_tmp_mut_46_sg1;
  reg [15:0] delta_conc_1_tmp_mut_47_sg1;
  reg [15:0] delta_conc_1_tmp_mut_48_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_49_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_50_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_51_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_52_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_53_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_54_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_55_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_56_sg1;
  reg [15:0] delta_conc_1_tmp_mut_49_sg1;
  reg [15:0] delta_conc_1_tmp_mut_50_sg1;
  reg [15:0] delta_conc_1_tmp_mut_51_sg1;
  reg [15:0] delta_conc_1_tmp_mut_52_sg1;
  reg [15:0] delta_conc_1_tmp_mut_53_sg1;
  reg [15:0] delta_conc_1_tmp_mut_54_sg1;
  reg [15:0] delta_conc_1_tmp_mut_55_sg1;
  reg [15:0] delta_conc_1_tmp_mut_56_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_57_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_58_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_59_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_60_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_61_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_62_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_63_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_64_sg1;
  reg [15:0] delta_conc_1_tmp_mut_57_sg1;
  reg [15:0] delta_conc_1_tmp_mut_58_sg1;
  reg [15:0] delta_conc_1_tmp_mut_59_sg1;
  reg [15:0] delta_conc_1_tmp_mut_60_sg1;
  reg [15:0] delta_conc_1_tmp_mut_61_sg1;
  reg [15:0] delta_conc_1_tmp_mut_62_sg1;
  reg [15:0] delta_conc_1_tmp_mut_63_sg1;
  reg [15:0] delta_conc_1_tmp_mut_64_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_65_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_66_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_67_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_68_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_69_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_70_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_71_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_72_sg1;
  reg [15:0] delta_conc_1_tmp_mut_65_sg1;
  reg [15:0] delta_conc_1_tmp_mut_66_sg1;
  reg [15:0] delta_conc_1_tmp_mut_67_sg1;
  reg [15:0] delta_conc_1_tmp_mut_68_sg1;
  reg [15:0] delta_conc_1_tmp_mut_69_sg1;
  reg [15:0] delta_conc_1_tmp_mut_70_sg1;
  reg [15:0] delta_conc_1_tmp_mut_71_sg1;
  reg [15:0] delta_conc_1_tmp_mut_72_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_73_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_74_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_75_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_76_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_77_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_78_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_79_sg1;
  reg [16:0] else_7_if_1_conc_tmp_mut_80_sg1;
  reg [15:0] delta_conc_1_tmp_mut_73_sg1;
  reg [15:0] delta_conc_1_tmp_mut_74_sg1;
  reg [15:0] delta_conc_1_tmp_mut_75_sg1;
  reg [15:0] delta_conc_1_tmp_mut_76_sg1;
  reg [15:0] delta_conc_1_tmp_mut_77_sg1;
  reg [15:0] delta_conc_1_tmp_mut_78_sg1;
  reg [15:0] delta_conc_1_tmp_mut_79_sg1;
  reg [15:0] delta_conc_1_tmp_mut_80_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_9_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_10_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_11_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_12_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_13_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_14_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_15_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_16_sg1;
  reg [15:0] max_conc_4_tmp_mut_9_sg1;
  reg [15:0] max_conc_4_tmp_mut_10_sg1;
  reg [15:0] max_conc_4_tmp_mut_11_sg1;
  reg [15:0] max_conc_4_tmp_mut_12_sg1;
  reg [15:0] max_conc_4_tmp_mut_13_sg1;
  reg [15:0] max_conc_4_tmp_mut_14_sg1;
  reg [15:0] max_conc_4_tmp_mut_15_sg1;
  reg [15:0] max_conc_4_tmp_mut_16_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_17_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_18_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_19_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_20_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_21_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_22_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_23_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_24_sg1;
  reg [15:0] max_conc_4_tmp_mut_17_sg1;
  reg [15:0] max_conc_4_tmp_mut_18_sg1;
  reg [15:0] max_conc_4_tmp_mut_19_sg1;
  reg [15:0] max_conc_4_tmp_mut_20_sg1;
  reg [15:0] max_conc_4_tmp_mut_21_sg1;
  reg [15:0] max_conc_4_tmp_mut_22_sg1;
  reg [15:0] max_conc_4_tmp_mut_23_sg1;
  reg [15:0] max_conc_4_tmp_mut_24_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_25_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_26_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_27_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_28_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_29_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_30_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_31_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_32_sg1;
  reg [15:0] max_conc_4_tmp_mut_25_sg1;
  reg [15:0] max_conc_4_tmp_mut_26_sg1;
  reg [15:0] max_conc_4_tmp_mut_27_sg1;
  reg [15:0] max_conc_4_tmp_mut_28_sg1;
  reg [15:0] max_conc_4_tmp_mut_29_sg1;
  reg [15:0] max_conc_4_tmp_mut_30_sg1;
  reg [15:0] max_conc_4_tmp_mut_31_sg1;
  reg [15:0] max_conc_4_tmp_mut_32_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_33_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_34_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_35_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_36_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_37_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_38_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_39_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_40_sg1;
  reg [15:0] max_conc_4_tmp_mut_33_sg1;
  reg [15:0] max_conc_4_tmp_mut_34_sg1;
  reg [15:0] max_conc_4_tmp_mut_35_sg1;
  reg [15:0] max_conc_4_tmp_mut_36_sg1;
  reg [15:0] max_conc_4_tmp_mut_37_sg1;
  reg [15:0] max_conc_4_tmp_mut_38_sg1;
  reg [15:0] max_conc_4_tmp_mut_39_sg1;
  reg [15:0] max_conc_4_tmp_mut_40_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_41_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_42_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_43_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_44_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_45_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_46_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_47_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_48_sg1;
  reg [15:0] max_conc_4_tmp_mut_41_sg1;
  reg [15:0] max_conc_4_tmp_mut_42_sg1;
  reg [15:0] max_conc_4_tmp_mut_43_sg1;
  reg [15:0] max_conc_4_tmp_mut_44_sg1;
  reg [15:0] max_conc_4_tmp_mut_45_sg1;
  reg [15:0] max_conc_4_tmp_mut_46_sg1;
  reg [15:0] max_conc_4_tmp_mut_47_sg1;
  reg [15:0] max_conc_4_tmp_mut_48_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_49_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_50_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_51_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_52_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_53_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_54_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_55_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_56_sg1;
  reg [15:0] max_conc_4_tmp_mut_49_sg1;
  reg [15:0] max_conc_4_tmp_mut_50_sg1;
  reg [15:0] max_conc_4_tmp_mut_51_sg1;
  reg [15:0] max_conc_4_tmp_mut_52_sg1;
  reg [15:0] max_conc_4_tmp_mut_53_sg1;
  reg [15:0] max_conc_4_tmp_mut_54_sg1;
  reg [15:0] max_conc_4_tmp_mut_55_sg1;
  reg [15:0] max_conc_4_tmp_mut_56_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_57_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_58_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_59_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_60_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_61_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_62_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_63_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_64_sg1;
  reg [15:0] max_conc_4_tmp_mut_57_sg1;
  reg [15:0] max_conc_4_tmp_mut_58_sg1;
  reg [15:0] max_conc_4_tmp_mut_59_sg1;
  reg [15:0] max_conc_4_tmp_mut_60_sg1;
  reg [15:0] max_conc_4_tmp_mut_61_sg1;
  reg [15:0] max_conc_4_tmp_mut_62_sg1;
  reg [15:0] max_conc_4_tmp_mut_63_sg1;
  reg [15:0] max_conc_4_tmp_mut_64_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_65_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_66_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_67_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_68_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_69_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_70_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_71_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_72_sg1;
  reg [15:0] max_conc_4_tmp_mut_65_sg1;
  reg [15:0] max_conc_4_tmp_mut_66_sg1;
  reg [15:0] max_conc_4_tmp_mut_67_sg1;
  reg [15:0] max_conc_4_tmp_mut_68_sg1;
  reg [15:0] max_conc_4_tmp_mut_69_sg1;
  reg [15:0] max_conc_4_tmp_mut_70_sg1;
  reg [15:0] max_conc_4_tmp_mut_71_sg1;
  reg [15:0] max_conc_4_tmp_mut_72_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_73_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_74_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_75_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_76_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_77_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_78_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_79_sg1;
  reg [15:0] else_7_if_conc_tmp_mut_80_sg1;
  reg [15:0] max_conc_4_tmp_mut_73_sg1;
  reg [15:0] max_conc_4_tmp_mut_74_sg1;
  reg [15:0] max_conc_4_tmp_mut_75_sg1;
  reg [15:0] max_conc_4_tmp_mut_76_sg1;
  reg [15:0] max_conc_4_tmp_mut_77_sg1;
  reg [15:0] max_conc_4_tmp_mut_78_sg1;
  reg [15:0] max_conc_4_tmp_mut_79_sg1;
  reg [15:0] max_conc_4_tmp_mut_80_sg1;
  wire and_506_cse;
  wire and_878_cse;
  wire and_1250_cse;
  wire and_1622_cse;
  wire and_1994_cse;
  wire and_2366_cse;
  wire and_2973_cse;
  wire and_2976_cse;
  wire and_2979_cse;
  wire and_2982_cse;
  wire and_2985_cse;
  wire and_2988_cse;
  wire and_2991_cse;
  wire and_2994_cse;
  wire and_2997_cse;
  wire and_3065_cse;
  wire and_3068_cse;
  wire and_3071_cse;
  wire and_3074_cse;
  wire and_3077_cse;
  wire and_3080_cse;
  wire and_3083_cse;
  wire and_3086_cse;
  wire and_3089_cse;
  wire [11:0] h_2_lpi_dfm_1_sg2_1;
  wire h_2_lpi_dfm_1_sg1_1;
  wire [16:0] h_2_lpi_dfm_4;
  wire or_303_cse;
  wire or_626_cse;
  wire or_628_cse;
  wire or_630_cse;
  wire and_3159_cse;
  wire and_3165_cse;
  wire or_605_cse;
  wire or_831_cse;
  wire or_833_cse;
  wire or_835_cse;
  wire and_3305_cse;
  wire or_1036_cse;
  wire or_1038_cse;
  wire or_1040_cse;
  wire and_3445_cse;
  wire or_1241_cse;
  wire or_1243_cse;
  wire or_1245_cse;
  wire and_3585_cse;
  wire or_1446_cse;
  wire or_1448_cse;
  wire or_1450_cse;
  wire and_3725_cse;
  wire or_1651_cse;
  wire or_1653_cse;
  wire or_1655_cse;
  wire and_3865_cse;
  wire or_1856_cse;
  wire or_1858_cse;
  wire or_1860_cse;
  wire and_4005_cse;
  wire or_2061_cse;
  wire nand_33_cse;
  wire or_2065_cse;
  wire and_4145_cse;
  wire or_2269_cse;
  wire or_2271_cse;
  wire or_2273_cse;
  wire and_4285_cse;
  wire mux_363_cse;
  wire mux_367_cse;
  wire and_4415_cse;
  wire and_4422_cse;
  wire and_4430_cse;
  wire mux_375_cse;
  wire mux_379_cse;
  wire and_4566_cse;
  wire and_4573_cse;
  wire and_4581_cse;
  wire mux_387_cse;
  wire mux_391_cse;
  wire and_4717_cse;
  wire and_4724_cse;
  wire and_4732_cse;
  wire mux_399_cse;
  wire mux_403_cse;
  wire and_4868_cse;
  wire and_4875_cse;
  wire and_4883_cse;
  wire mux_411_cse;
  wire mux_415_cse;
  wire and_5019_cse;
  wire and_5026_cse;
  wire and_5034_cse;
  wire mux_423_cse;
  wire mux_427_cse;
  wire and_5170_cse;
  wire and_5177_cse;
  wire and_5185_cse;
  wire mux_435_cse;
  wire mux_439_cse;
  wire and_5321_cse;
  wire and_5328_cse;
  wire and_5336_cse;
  wire mux_447_cse;
  wire mux_451_cse;
  wire and_5472_cse;
  wire and_5479_cse;
  wire and_5487_cse;
  wire and_5623_cse;
  wire and_5630_cse;
  wire and_5638_cse;
  wire and_5737_cse;
  wire and_5745_cse;
  wire and_5754_cse;
  wire and_5763_cse;
  wire and_5904_cse;
  wire and_5912_cse;
  wire and_5921_cse;
  wire and_5930_cse;
  wire and_6071_cse;
  wire and_6079_cse;
  wire and_6088_cse;
  wire and_6097_cse;
  wire and_6238_cse;
  wire and_6246_cse;
  wire and_6255_cse;
  wire and_6264_cse;
  wire and_6405_cse;
  wire and_6413_cse;
  wire and_6422_cse;
  wire and_6431_cse;
  wire and_6572_cse;
  wire and_6580_cse;
  wire and_6589_cse;
  wire and_6598_cse;
  wire and_6739_cse;
  wire and_6747_cse;
  wire and_6756_cse;
  wire and_6765_cse;
  wire and_6906_cse;
  wire and_6914_cse;
  wire and_6923_cse;
  wire and_6932_cse;
  wire and_7073_cse;
  wire and_7081_cse;
  wire and_7090_cse;
  wire and_7204_cse;
  wire and_7212_cse;
  wire and_7221_cse;
  wire and_7231_cse;
  wire and_7242_cse;
  wire and_7254_cse;
  wire and_7267_cse;
  wire and_7281_cse;
  wire and_7288_cse;
  wire and_7383_cse;
  wire and_7391_cse;
  wire and_7400_cse;
  wire and_7410_cse;
  wire and_7421_cse;
  wire and_7433_cse;
  wire and_7446_cse;
  wire and_7460_cse;
  wire and_7467_cse;
  wire and_7562_cse;
  wire and_7570_cse;
  wire and_7579_cse;
  wire and_7589_cse;
  wire and_7600_cse;
  wire and_7612_cse;
  wire and_7625_cse;
  wire and_7639_cse;
  wire and_7646_cse;
  wire and_7741_cse;
  wire and_7749_cse;
  wire and_7758_cse;
  wire and_7768_cse;
  wire and_7779_cse;
  wire and_7791_cse;
  wire and_7804_cse;
  wire and_7818_cse;
  wire and_7825_cse;
  wire and_7920_cse;
  wire and_7928_cse;
  wire and_7937_cse;
  wire and_7947_cse;
  wire and_7958_cse;
  wire and_7970_cse;
  wire and_7983_cse;
  wire and_7997_cse;
  wire and_8004_cse;
  wire and_8099_cse;
  wire and_8107_cse;
  wire and_8116_cse;
  wire and_8126_cse;
  wire and_8137_cse;
  wire and_8149_cse;
  wire and_8162_cse;
  wire and_8176_cse;
  wire and_8183_cse;
  wire and_8278_cse;
  wire and_8286_cse;
  wire and_8295_cse;
  wire and_8305_cse;
  wire and_8316_cse;
  wire and_8328_cse;
  wire and_8341_cse;
  wire and_8355_cse;
  wire and_8362_cse;
  wire and_8457_cse;
  wire and_8465_cse;
  wire and_8474_cse;
  wire and_8484_cse;
  wire and_8495_cse;
  wire and_8507_cse;
  wire and_8520_cse;
  wire and_8534_cse;
  wire and_8541_cse;
  wire and_8636_cse;
  wire and_8644_cse;
  wire and_8653_cse;
  wire and_8663_cse;
  wire and_9058_cse;
  wire and_2924_cse;
  wire and_3062_cse;
  wire and_3154_cse;
  wire or_5023_cse;
  wire or_5033_cse;
  wire or_5043_cse;
  wire or_5053_cse;
  wire or_5063_cse;
  wire or_5073_cse;
  wire or_5083_cse;
  wire or_5093_cse;
  wire or_5103_cse;
  wire or_5114_cse;
  wire or_5126_cse;
  wire or_5138_cse;
  wire or_5150_cse;
  wire or_5162_cse;
  wire or_5174_cse;
  wire or_5186_cse;
  wire or_5198_cse;
  wire or_5210_cse;
  wire or_5222_cse;
  wire or_5234_cse;
  wire or_5246_cse;
  wire or_5258_cse;
  wire or_5270_cse;
  wire or_5282_cse;
  wire or_5294_cse;
  wire or_5306_cse;
  wire or_5318_cse;
  wire or_612_cse;
  wire or_817_cse;
  wire or_1022_cse;
  wire or_1227_cse;
  wire or_1432_cse;
  wire or_1637_cse;
  wire or_1842_cse;
  wire nand_cse;
  wire or_2252_cse;
  reg [15:0] reg_div_mgc_div_28_b_tmp;
  reg [15:0] reg_div_mgc_div_28_a_tmp;
  reg [15:0] reg_div_mgc_div_29_b_tmp;
  reg [15:0] reg_div_mgc_div_29_a_tmp;
  reg [15:0] reg_div_mgc_div_30_b_tmp;
  reg [15:0] reg_div_mgc_div_30_a_tmp;
  reg [15:0] reg_div_mgc_div_31_b_tmp;
  reg [15:0] reg_div_mgc_div_31_a_tmp;
  reg [15:0] reg_div_mgc_div_32_b_tmp;
  reg [15:0] reg_div_mgc_div_32_a_tmp;
  reg [15:0] reg_div_mgc_div_33_b_tmp;
  reg [15:0] reg_div_mgc_div_33_a_tmp;
  reg [15:0] reg_div_mgc_div_34_b_tmp;
  reg [15:0] reg_div_mgc_div_34_a_tmp;
  reg [15:0] reg_div_mgc_div_35_b_tmp;
  reg [15:0] reg_div_mgc_div_35_a_tmp;
  reg [15:0] reg_div_mgc_div_27_b_tmp;
  reg [15:0] reg_div_mgc_div_27_a_tmp;
  reg [15:0] reg_div_mgc_div_19_b_tmp;
  reg [16:0] reg_div_mgc_div_19_a_tmp;
  reg [15:0] reg_div_mgc_div_20_b_tmp;
  reg [16:0] reg_div_mgc_div_20_a_tmp;
  reg [15:0] reg_div_mgc_div_21_b_tmp;
  reg [16:0] reg_div_mgc_div_21_a_tmp;
  reg [15:0] reg_div_mgc_div_22_b_tmp;
  reg [16:0] reg_div_mgc_div_22_a_tmp;
  reg [15:0] reg_div_mgc_div_23_b_tmp;
  reg [16:0] reg_div_mgc_div_23_a_tmp;
  reg [15:0] reg_div_mgc_div_24_b_tmp;
  reg [16:0] reg_div_mgc_div_24_a_tmp;
  reg [15:0] reg_div_mgc_div_25_b_tmp;
  reg [16:0] reg_div_mgc_div_25_a_tmp;
  reg [15:0] reg_div_mgc_div_26_b_tmp;
  reg [16:0] reg_div_mgc_div_26_a_tmp;
  reg [15:0] reg_div_mgc_div_b_tmp;
  reg [16:0] reg_div_mgc_div_a_tmp;
  reg [15:0] reg_div_mgc_div_10_b_tmp;
  reg [16:0] reg_div_mgc_div_10_a_tmp;
  reg [15:0] reg_div_mgc_div_11_b_tmp;
  reg [16:0] reg_div_mgc_div_11_a_tmp;
  reg [15:0] reg_div_mgc_div_12_b_tmp;
  reg [16:0] reg_div_mgc_div_12_a_tmp;
  reg [15:0] reg_div_mgc_div_13_b_tmp;
  reg [16:0] reg_div_mgc_div_13_a_tmp;
  reg [15:0] reg_div_mgc_div_14_b_tmp;
  reg [16:0] reg_div_mgc_div_14_a_tmp;
  reg [15:0] reg_div_mgc_div_15_b_tmp;
  reg [16:0] reg_div_mgc_div_15_a_tmp;
  reg [15:0] reg_div_mgc_div_16_b_tmp;
  reg [16:0] reg_div_mgc_div_16_a_tmp;
  reg [15:0] reg_div_mgc_div_17_b_tmp;
  reg [16:0] reg_div_mgc_div_17_a_tmp;
  reg [15:0] reg_div_mgc_div_18_b_tmp;
  reg [16:0] reg_div_mgc_div_18_a_tmp;
  reg [15:0] reg_div_mgc_div_1_b_tmp;
  reg [16:0] reg_div_mgc_div_1_a_tmp;
  reg [15:0] reg_div_mgc_div_2_b_tmp;
  reg [16:0] reg_div_mgc_div_2_a_tmp;
  reg [15:0] reg_div_mgc_div_3_b_tmp;
  reg [16:0] reg_div_mgc_div_3_a_tmp;
  reg [15:0] reg_div_mgc_div_4_b_tmp;
  reg [16:0] reg_div_mgc_div_4_a_tmp;
  reg [15:0] reg_div_mgc_div_5_b_tmp;
  reg [16:0] reg_div_mgc_div_5_a_tmp;
  reg [15:0] reg_div_mgc_div_6_b_tmp;
  reg [16:0] reg_div_mgc_div_6_a_tmp;
  reg [15:0] reg_div_mgc_div_7_b_tmp;
  reg [16:0] reg_div_mgc_div_7_a_tmp;
  reg [15:0] reg_div_mgc_div_8_b_tmp;
  reg [16:0] reg_div_mgc_div_8_a_tmp;
  reg [15:0] reg_div_mgc_div_9_b_tmp;
  reg [16:0] reg_div_mgc_div_9_a_tmp;
  wire mux_95_cse;
  wire mux_124_cse;
  wire and_3299_cse;
  wire mux_153_cse;
  wire and_3439_cse;
  wire mux_182_cse;
  wire and_3579_cse;
  wire mux_213_cse;
  wire and_3719_cse;
  wire mux_242_cse;
  wire and_3859_cse;
  wire mux_271_cse;
  wire and_3999_cse;
  wire and_4139_cse;
  wire mux_333_cse;
  wire and_4279_cse;
  wire and_4438_cse;
  wire and_4447_cse;
  wire and_4457_cse;
  wire and_4468_cse;
  wire and_4480_cse;
  wire and_4486_cse;
  wire and_4589_cse;
  wire and_4598_cse;
  wire and_4608_cse;
  wire and_4619_cse;
  wire and_4631_cse;
  wire and_4637_cse;
  wire and_4740_cse;
  wire and_4749_cse;
  wire and_4759_cse;
  wire and_4770_cse;
  wire and_4782_cse;
  wire and_4788_cse;
  wire and_4891_cse;
  wire and_4900_cse;
  wire and_4910_cse;
  wire and_4921_cse;
  wire and_4933_cse;
  wire and_4939_cse;
  wire and_5042_cse;
  wire and_5051_cse;
  wire and_5061_cse;
  wire and_5072_cse;
  wire and_5084_cse;
  wire and_5090_cse;
  wire and_5193_cse;
  wire and_5202_cse;
  wire and_5212_cse;
  wire and_5223_cse;
  wire and_5235_cse;
  wire and_5241_cse;
  wire and_5344_cse;
  wire and_5353_cse;
  wire and_5363_cse;
  wire and_5374_cse;
  wire and_5386_cse;
  wire and_5392_cse;
  wire and_5495_cse;
  wire and_5504_cse;
  wire and_5514_cse;
  wire and_5525_cse;
  wire and_5537_cse;
  wire and_5543_cse;
  wire and_5645_cse;
  wire and_5773_cse;
  wire and_5784_cse;
  wire and_5796_cse;
  wire and_5809_cse;
  wire mux_514_cse;
  wire and_5940_cse;
  wire and_5951_cse;
  wire and_5963_cse;
  wire and_5976_cse;
  wire mux_526_cse;
  wire and_6107_cse;
  wire and_6118_cse;
  wire and_6130_cse;
  wire and_6143_cse;
  wire mux_538_cse;
  wire and_6274_cse;
  wire and_6285_cse;
  wire and_6297_cse;
  wire and_6310_cse;
  wire mux_550_cse;
  wire and_6441_cse;
  wire and_6452_cse;
  wire and_6464_cse;
  wire and_6477_cse;
  wire mux_562_cse;
  wire and_6608_cse;
  wire and_6619_cse;
  wire and_6631_cse;
  wire and_6644_cse;
  wire mux_574_cse;
  wire and_6775_cse;
  wire and_6786_cse;
  wire and_6798_cse;
  wire and_6811_cse;
  wire mux_586_cse;
  wire and_6942_cse;
  wire and_6953_cse;
  wire and_6965_cse;
  wire and_6978_cse;
  wire mux_598_cse;
  wire and_7099_cse;
  wire and_8673_cse;
  wire or_4933_cse;
  wire or_4943_cse;
  wire or_4953_cse;
  wire or_4963_cse;
  wire or_4973_cse;
  wire or_4983_cse;
  wire or_4993_cse;
  wire or_5003_cse;
  wire or_5013_cse;
  wire or_5325_cse;
  wire mux_460_cse;
  wire and_2362_cse;
  wire and_1990_cse;
  wire and_1618_cse;
  wire and_1246_cse;
  wire and_874_cse;
  wire and_502_cse;
  wire and_9092_cse;
  wire and_3207_cse;
  wire and_3347_cse;
  wire and_3487_cse;
  wire and_3627_cse;
  wire and_3767_cse;
  wire and_3907_cse;
  wire and_4047_cse;
  wire mux_302_cse;
  wire and_4195_cse;
  wire and_4325_cse;
  wire mux_466_cse;
  wire mux_610_cse;
  wire mux_659_cse;
  wire and_3172_cse;
  wire and_3180_cse;
  wire and_3189_cse;
  wire and_3199_cse;
  wire and_3221_cse;
  wire and_3312_cse;
  wire and_3320_cse;
  wire and_3329_cse;
  wire and_3339_cse;
  wire and_3361_cse;
  wire and_3452_cse;
  wire and_3460_cse;
  wire and_3469_cse;
  wire and_3479_cse;
  wire and_3501_cse;
  wire and_3592_cse;
  wire and_3600_cse;
  wire and_3609_cse;
  wire and_3619_cse;
  wire and_3641_cse;
  wire and_3732_cse;
  wire and_3740_cse;
  wire and_3749_cse;
  wire and_3759_cse;
  wire and_3781_cse;
  wire and_3872_cse;
  wire and_3880_cse;
  wire and_3889_cse;
  wire and_3899_cse;
  wire and_3921_cse;
  wire and_4012_cse;
  wire and_4020_cse;
  wire and_4029_cse;
  wire and_4039_cse;
  wire and_4061_cse;
  wire and_4152_cse;
  wire and_4160_cse;
  wire and_4291_cse;
  wire and_4298_cse;
  wire and_4307_cse;
  wire and_4317_cse;
  wire and_4339_cse;
  wire and_7108_cse;
  wire and_4187_cse;
  wire mux_471_cse;
  wire mux_615_cse;
  wire mux_664_cse;
  wire and_8701_cse;
  wire and_3209_cse;
  wire and_3349_cse;
  wire and_3489_cse;
  wire and_3629_cse;
  wire and_3769_cse;
  wire and_3909_cse;
  wire and_4049_cse;
  wire and_4169_cse;
  wire and_4179_cse;
  wire and_4201_cse;
  wire and_4327_cse;
  wire and_5652_cse;
  wire and_7116_cse;
  wire and_8682_cse;
  wire mux_105_cse;
  wire mux_134_cse;
  wire mux_163_cse;
  wire mux_192_cse;
  wire mux_223_cse;
  wire mux_252_cse;
  wire mux_281_cse;
  wire mux_343_cse;
  wire mux_476_cse;
  wire mux_621_cse;
  wire mux_627_cse;
  wire and_4189_cse;
  wire and_5659_cse;
  wire and_5666_cse;
  wire and_7124_cse;
  wire and_8691_cse;
  wire and_8700_cse;
  wire and_8702_cse;
  wire mux_310_cse;
  wire mux_482_cse;
  wire mux_106_cse;
  wire mux_135_cse;
  wire mux_164_cse;
  wire mux_194_cse;
  wire mux_224_cse;
  wire mux_253_cse;
  wire mux_282_cse;
  wire mux_345_cse;
  wire and_7132_cse;
  wire mux_628_cse;
  wire mux_312_cse;
  wire and_5674_cse;
  wire mux_483_cse;
  wire [29:0] else_7_acc_2_itm;
  wire [30:0] nl_else_7_acc_2_itm;
  wire [15:0] else_7_acc_2_psp_sg1_sva_1;
  wire [29:0] h_2_sva_duc_mx0;
  wire [12:0] h_2_sva_1_sg1;
  wire [13:0] nl_h_2_sva_1_sg1;
  wire [29:0] div_sdt_3_sva_duc_mx0;
  wire else_7_nor_ssc;
  wire [3:0] else_7_if_acc_idiv;
  wire [4:0] nl_else_7_if_acc_idiv;
  wire [3:0] else_7_if_1_acc_idiv;
  wire [4:0] nl_else_7_if_1_acc_idiv;
  wire [15:0] g_sg1_lpi_dfm;
  wire [15:0] b_sg1_lpi_dfm;
  wire [3:0] else_7_else_1_if_acc_idiv;
  wire [4:0] nl_else_7_else_1_if_acc_idiv;
  wire [15:0] r_sg1_lpi_dfm;
  wire [3:0] else_7_else_1_else_acc_idiv;
  wire [4:0] nl_else_7_else_1_else_acc_idiv;
  wire unequal_tmp;
  wire [15:0] min_sg1_lpi_dfm_3;
  wire [17:0] if_if_acc_1_itm;
  wire [18:0] nl_if_if_acc_1_itm;
  wire [17:0] else_1_if_acc_1_itm;
  wire [18:0] nl_else_1_if_acc_1_itm;
  wire [17:0] if_3_if_acc_1_itm;
  wire [18:0] nl_if_3_if_acc_1_itm;
  wire [17:0] else_5_if_acc_1_itm;
  wire [18:0] nl_else_5_if_acc_1_itm;
  wire [16:0] else_7_acc_3_itm;
  wire [17:0] nl_else_7_acc_3_itm;
  wire [4:0] acc_5_itm;
  wire [5:0] nl_acc_5_itm;
  wire [17:0] else_7_if_1_acc_1_itm;
  wire [18:0] nl_else_7_if_1_acc_1_itm;
  wire [4:0] acc_itm;
  wire [5:0] nl_acc_itm;
  wire [17:0] else_7_else_1_if_acc_2_itm;
  wire [18:0] nl_else_7_else_1_if_acc_2_itm;
  wire [4:0] acc_6_itm;
  wire [5:0] nl_acc_6_itm;
  wire [17:0] else_7_else_1_else_acc_2_itm;
  wire [18:0] nl_else_7_else_1_else_acc_2_itm;
  wire [4:0] acc_7_itm;
  wire [5:0] nl_acc_7_itm;
  wire [17:0] if_3_acc_itm;
  wire [18:0] nl_if_3_acc_itm;
  wire [17:0] if_acc_itm;
  wire [18:0] nl_if_acc_itm;

  wire[0:0] mux_92_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] mux_653_nl;
  wire[12:0] mux1h_5_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] mux_670_nl;

  // Interconnect Declarations for Component Instantiations 
  assign or_303_cse = (max_sg1_lpi_dfm_3_st_9[15]) | (max_sg1_lpi_dfm_3_st_9[14])
      | (max_sg1_lpi_dfm_3_st_9[13]) | (max_sg1_lpi_dfm_3_st_9[12]) | (max_sg1_lpi_dfm_3_st_9[11])
      | (max_sg1_lpi_dfm_3_st_9[10]) | (max_sg1_lpi_dfm_3_st_9[9]) | (max_sg1_lpi_dfm_3_st_9[8])
      | (max_sg1_lpi_dfm_3_st_9[7]) | (max_sg1_lpi_dfm_3_st_9[6]) | (max_sg1_lpi_dfm_3_st_9[5])
      | (max_sg1_lpi_dfm_3_st_9[4]) | (max_sg1_lpi_dfm_3_st_9[3]) | (max_sg1_lpi_dfm_3_st_9[2])
      | (max_sg1_lpi_dfm_3_st_9[1]) | (max_sg1_lpi_dfm_3_st_9[0]);
  assign and_9092_cse = (~ if_7_equal_svs_9) & main_stage_0_10;
  assign and_2924_cse = ((else_7_if_1_div_9cyc_st_9[0]) | (else_7_if_1_div_9cyc_st_9[1])
      | (else_7_if_1_div_9cyc_st_9[2])) & (else_7_if_1_div_9cyc_st_9[3]);
  assign and_3062_cse = ((else_7_else_1_if_div_9cyc_st_9[2]) | (else_7_else_1_if_div_9cyc_st_9[1])
      | (else_7_else_1_if_div_9cyc_st_9[0])) & (else_7_else_1_if_div_9cyc_st_9[3]);
  assign and_3154_cse = ((else_7_else_1_else_div_9cyc_st_9[0]) | (else_7_else_1_else_div_9cyc_st_9[1])
      | (else_7_else_1_else_div_9cyc_st_9[2])) & (else_7_else_1_else_div_9cyc_st_9[3]);
  assign or_626_cse = (~ or_tmp_7) | (else_7_if_acc_tmp[0]) | (else_7_if_acc_tmp[1])
      | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign or_628_cse = (~ or_tmp_6) | (else_7_if_div_9cyc_st_1[0]) | (else_7_if_div_9cyc_st_1[1])
      | (else_7_if_div_9cyc_st_1[2]) | (else_7_if_div_9cyc_st_1[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_630_cse = (~ or_tmp_28) | (else_7_if_div_9cyc_st_2[2]) | (else_7_if_div_9cyc_st_2[1])
      | (else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign or_605_cse = (mux1h_81_tmp[0]) | (mux1h_81_tmp[1]) | (mux1h_81_tmp[2]) |
      (mux1h_81_tmp[3]) | (mux1h_81_tmp[4]) | (mux1h_81_tmp[5]) | (mux1h_81_tmp[6])
      | (mux1h_81_tmp[7]) | (mux1h_81_tmp[8]) | (mux1h_81_tmp[9]) | (mux1h_81_tmp[10])
      | (mux1h_81_tmp[11]) | (mux1h_81_tmp[12]) | (mux1h_81_tmp[13]) | (mux1h_81_tmp[14])
      | (mux1h_81_tmp[15]);
  assign and_3159_cse = or_605_cse & and_dcpl_3146 & and_dcpl_3144;
  assign mux_92_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (else_7_if_acc_tmp[0])
      | (else_7_if_acc_tmp[1]) | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_3165_cse = (mux_92_nl) & and_dcpl_3152 & and_dcpl_3150;
  assign mux_95_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_31))) , or_tmp_31},
      or_630_cse);
  assign div_mgc_div_28_b = {reg_div_mgc_div_28_b_tmp , 16'b0};
  assign div_mgc_div_28_a = {reg_div_mgc_div_28_a_tmp , 32'b0};
  assign or_831_cse = (~ or_tmp_7) | (~ (else_7_if_acc_tmp[0])) | (else_7_if_acc_tmp[1])
      | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign or_833_cse = (~ or_tmp_6) | (~ (else_7_if_div_9cyc_st_1[0])) | (else_7_if_div_9cyc_st_1[1])
      | (else_7_if_div_9cyc_st_1[2]) | (else_7_if_div_9cyc_st_1[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_835_cse = (~ or_tmp_28) | (else_7_if_div_9cyc_st_2[2]) | (else_7_if_div_9cyc_st_2[1])
      | (~ (else_7_if_div_9cyc_st_2[0])) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign mux_121_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (~ (else_7_if_acc_tmp[0]))
      | (else_7_if_acc_tmp[1]) | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_3305_cse = (mux_121_nl) & and_dcpl_3152 & and_dcpl_3149 & (else_7_if_div_9cyc_st_1[0]);
  assign and_3299_cse = or_605_cse & and_dcpl_3146 & and_dcpl_3238;
  assign mux_124_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_206))) , or_tmp_206},
      or_835_cse);
  assign div_mgc_div_29_b = {reg_div_mgc_div_29_b_tmp , 16'b0};
  assign div_mgc_div_29_a = {reg_div_mgc_div_29_a_tmp , 32'b0};
  assign or_1036_cse = (~ or_tmp_7) | (else_7_if_acc_tmp[0]) | (~ (else_7_if_acc_tmp[1]))
      | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign or_1038_cse = (~ or_tmp_6) | (else_7_if_div_9cyc_st_1[0]) | (~ (else_7_if_div_9cyc_st_1[1]))
      | (else_7_if_div_9cyc_st_1[2]) | (else_7_if_div_9cyc_st_1[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_1040_cse = (~ or_tmp_28) | (else_7_if_div_9cyc_st_2[2]) | (~ (else_7_if_div_9cyc_st_2[1]))
      | (else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign mux_150_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (else_7_if_acc_tmp[0])
      | (~ (else_7_if_acc_tmp[1])) | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_3445_cse = (mux_150_nl) & and_dcpl_3152 & and_dcpl_3337 & (~ (else_7_if_div_9cyc_st_1[0]));
  assign and_3439_cse = or_605_cse & and_dcpl_3146 & and_dcpl_3332;
  assign mux_153_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_381))) , or_tmp_381},
      or_1040_cse);
  assign div_mgc_div_30_b = {reg_div_mgc_div_30_b_tmp , 16'b0};
  assign div_mgc_div_30_a = {reg_div_mgc_div_30_a_tmp , 32'b0};
  assign or_1241_cse = (~ or_tmp_7) | (~ (else_7_if_acc_tmp[0])) | (~ (else_7_if_acc_tmp[1]))
      | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign or_1243_cse = (~ or_tmp_6) | (~ (else_7_if_div_9cyc_st_1[0])) | (~ (else_7_if_div_9cyc_st_1[1]))
      | (else_7_if_div_9cyc_st_1[2]) | (else_7_if_div_9cyc_st_1[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_1245_cse = (~ or_tmp_28) | (else_7_if_div_9cyc_st_2[2]) | (~ (else_7_if_div_9cyc_st_2[1]))
      | (~ (else_7_if_div_9cyc_st_2[0])) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign mux_179_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (~ (else_7_if_acc_tmp[0]))
      | (~ (else_7_if_acc_tmp[1])) | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_3585_cse = (mux_179_nl) & and_dcpl_3152 & and_dcpl_3337 & (else_7_if_div_9cyc_st_1[0]);
  assign and_3579_cse = or_605_cse & and_dcpl_3146 & and_dcpl_3426;
  assign mux_182_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_556))) , or_tmp_556},
      or_1245_cse);
  assign div_mgc_div_31_b = {reg_div_mgc_div_31_b_tmp , 16'b0};
  assign div_mgc_div_31_a = {reg_div_mgc_div_31_a_tmp , 32'b0};
  assign or_1446_cse = (~ or_tmp_7) | (else_7_if_acc_tmp[0]) | (else_7_if_acc_tmp[1])
      | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign or_1448_cse = (~ or_tmp_6) | (else_7_if_div_9cyc_st_1[0]) | (else_7_if_div_9cyc_st_1[1])
      | (~ (else_7_if_div_9cyc_st_1[2])) | (else_7_if_div_9cyc_st_1[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_1450_cse = (~ or_tmp_28) | (~ (else_7_if_div_9cyc_st_2[2])) | (else_7_if_div_9cyc_st_2[1])
      | (else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign mux_210_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (else_7_if_acc_tmp[0])
      | (else_7_if_acc_tmp[1]) | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_3725_cse = (mux_210_nl) & and_dcpl_3152 & and_dcpl_3525 & (~ (else_7_if_div_9cyc_st_1[0]));
  assign and_3719_cse = or_605_cse & and_dcpl_3522 & and_dcpl_3144;
  assign mux_213_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_731))) , or_tmp_731},
      or_1450_cse);
  assign div_mgc_div_32_b = {reg_div_mgc_div_32_b_tmp , 16'b0};
  assign div_mgc_div_32_a = {reg_div_mgc_div_32_a_tmp , 32'b0};
  assign or_1651_cse = (~ or_tmp_7) | (~ (else_7_if_acc_tmp[0])) | (else_7_if_acc_tmp[1])
      | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign or_1653_cse = (~ or_tmp_6) | (~ (else_7_if_div_9cyc_st_1[0])) | (else_7_if_div_9cyc_st_1[1])
      | (~ (else_7_if_div_9cyc_st_1[2])) | (else_7_if_div_9cyc_st_1[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_1655_cse = (~ or_tmp_28) | (~ (else_7_if_div_9cyc_st_2[2])) | (else_7_if_div_9cyc_st_2[1])
      | (~ (else_7_if_div_9cyc_st_2[0])) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign mux_239_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (~ (else_7_if_acc_tmp[0]))
      | (else_7_if_acc_tmp[1]) | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_3865_cse = (mux_239_nl) & and_dcpl_3152 & and_dcpl_3525 & (else_7_if_div_9cyc_st_1[0]);
  assign and_3859_cse = or_605_cse & and_dcpl_3522 & and_dcpl_3238;
  assign mux_242_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_906))) , or_tmp_906},
      or_1655_cse);
  assign div_mgc_div_33_b = {reg_div_mgc_div_33_b_tmp , 16'b0};
  assign div_mgc_div_33_a = {reg_div_mgc_div_33_a_tmp , 32'b0};
  assign or_1856_cse = (~ or_tmp_7) | (else_7_if_acc_tmp[0]) | (~ (else_7_if_acc_tmp[1]))
      | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign or_1858_cse = (~ or_tmp_6) | (else_7_if_div_9cyc_st_1[0]) | (~ (else_7_if_div_9cyc_st_1[1]))
      | (~ (else_7_if_div_9cyc_st_1[2])) | (else_7_if_div_9cyc_st_1[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_1860_cse = (~ or_tmp_28) | (~ (else_7_if_div_9cyc_st_2[2])) | (~ (else_7_if_div_9cyc_st_2[1]))
      | (else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign mux_268_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (else_7_if_acc_tmp[0])
      | (~ (else_7_if_acc_tmp[1])) | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_4005_cse = (mux_268_nl) & and_dcpl_3152 & and_dcpl_3713 & (~ (else_7_if_div_9cyc_st_1[0]));
  assign and_3999_cse = or_605_cse & and_dcpl_3522 & and_dcpl_3332;
  assign mux_271_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_1081))) , or_tmp_1081},
      or_1860_cse);
  assign div_mgc_div_34_b = {reg_div_mgc_div_34_b_tmp , 16'b0};
  assign div_mgc_div_34_a = {reg_div_mgc_div_34_a_tmp , 32'b0};
  assign or_2061_cse = (~ or_tmp_7) | (~ (else_7_if_acc_tmp[0])) | (~ (else_7_if_acc_tmp[1]))
      | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3]) | if_7_equal_tmp;
  assign nand_33_cse = ~(or_tmp_6 & (else_7_if_div_9cyc_st_1[0]) & (else_7_if_div_9cyc_st_1[1])
      & (else_7_if_div_9cyc_st_1[2]) & (~ (else_7_if_div_9cyc_st_1[3])) & main_stage_0_2
      & (~ if_7_equal_svs_st_1));
  assign or_2065_cse = (~ or_tmp_28) | (~ (else_7_if_div_9cyc_st_2[2])) | (~ (else_7_if_div_9cyc_st_2[1]))
      | (~ (else_7_if_div_9cyc_st_2[0])) | (else_7_if_div_9cyc_st_2[3]) | if_7_equal_svs_st_2;
  assign mux_297_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (~ (else_7_if_acc_tmp[0]))
      | (~ (else_7_if_acc_tmp[1])) | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[3])
      | if_7_equal_tmp);
  assign and_4145_cse = (mux_297_nl) & and_dcpl_3152 & and_dcpl_3713 & (else_7_if_div_9cyc_st_1[0]);
  assign and_4139_cse = or_605_cse & and_dcpl_3522 & and_dcpl_3426;
  assign div_mgc_div_35_b = {reg_div_mgc_div_35_b_tmp , 16'b0};
  assign div_mgc_div_35_a = {reg_div_mgc_div_35_a_tmp , 32'b0};
  assign or_2269_cse = (~ or_tmp_7) | (else_7_if_acc_tmp[0]) | (else_7_if_acc_tmp[1])
      | (else_7_if_acc_tmp[2]) | (~ (else_7_if_acc_tmp[3])) | if_7_equal_tmp;
  assign or_2271_cse = (~ or_tmp_6) | (else_7_if_div_9cyc_st_1[0]) | (else_7_if_div_9cyc_st_1[1])
      | (else_7_if_div_9cyc_st_1[2]) | (~ (else_7_if_div_9cyc_st_1[3])) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_2273_cse = (~ or_tmp_28) | (else_7_if_div_9cyc_st_2[2]) | (else_7_if_div_9cyc_st_2[1])
      | (else_7_if_div_9cyc_st_2[0]) | (~ (else_7_if_div_9cyc_st_2[3])) | if_7_equal_svs_st_2;
  assign mux_328_nl = MUX_s_1_2_2({not_tmp_146 , or_tmp_6}, (else_7_if_acc_tmp[0])
      | (else_7_if_acc_tmp[1]) | (else_7_if_acc_tmp[2]) | (~ (else_7_if_acc_tmp[3]))
      | if_7_equal_tmp);
  assign and_4285_cse = (mux_328_nl) & and_2366_cse & (else_7_if_div_9cyc_st_1[3])
      & and_dcpl_3150;
  assign and_4279_cse = or_605_cse & (~ if_7_equal_tmp) & (else_7_if_acc_tmp[3])
      & (~ (else_7_if_acc_tmp[2])) & and_dcpl_3144;
  assign mux_333_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_1434))) , or_tmp_1434},
      or_2273_cse);
  assign div_mgc_div_27_b = {reg_div_mgc_div_27_b_tmp , 16'b0};
  assign div_mgc_div_27_a = {reg_div_mgc_div_27_a_tmp , 32'b0};
  assign mux_363_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_1593)))
      , or_tmp_1593}, or_tmp_1592);
  assign mux_367_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_421)))
      , and_tmp_421}, or_tmp_1592);
  assign and_4415_cse = and_dcpl_3993 & and_dcpl_3991;
  assign and_4422_cse = (~((~(or_dcpl_857 | or_dcpl_855)) | if_7_equal_svs_st_1))
      & and_dcpl_3998 & and_dcpl_3996;
  assign and_4430_cse = ((else_7_if_1_acc_tmp[2]) | (else_7_if_1_acc_tmp[0]) | (else_7_if_1_acc_tmp[3])
      | (else_7_if_1_acc_tmp[1]) | (~ else_7_equal_tmp) | if_7_equal_tmp) & ((else_7_if_1_div_9cyc[0])
      | (else_7_if_1_div_9cyc[1]) | (else_7_if_1_div_9cyc[3]) | (else_7_if_1_div_9cyc[2])
      | (~ else_7_equal_svs_st_1) | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4006
      & and_dcpl_4003;
  assign and_4438_cse = or_tmp_1591 & mux_363_cse & and_dcpl_4013 & and_dcpl_4010;
  assign and_4447_cse = or_tmp_1595 & or_tmp_1591 & mux_363_cse & and_dcpl_4020 &
      and_dcpl_4017;
  assign and_4457_cse = or_tmp_1600 & or_tmp_1595 & or_tmp_1591 & mux_363_cse & and_dcpl_4027
      & and_dcpl_4024;
  assign and_4468_cse = or_tmp_1606 & or_tmp_1600 & or_tmp_1595 & or_tmp_1591 & mux_363_cse
      & and_dcpl_4034 & and_dcpl_4031;
  assign and_4480_cse = or_tmp_1613 & or_tmp_1606 & or_tmp_1600 & or_tmp_1595 & mux_367_cse
      & and_dcpl_4041 & and_dcpl_4038;
  assign and_4486_cse = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (else_7_if_1_div_9cyc_st_7[0]) | (else_7_if_1_div_9cyc_st_7[1]) | (else_7_if_1_div_9cyc_st_7[2])
      | (else_7_if_1_div_9cyc_st_7[3])) & or_tmp_1613 & or_tmp_1606 & or_tmp_1600
      & or_tmp_1595 & mux_367_cse;
  assign div_mgc_div_19_b = {reg_div_mgc_div_19_b_tmp , 16'b0};
  assign div_mgc_div_19_a = {reg_div_mgc_div_19_a_tmp , 32'b0};
  assign mux_375_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_1673)))
      , or_tmp_1673}, or_tmp_1672);
  assign mux_379_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_464)))
      , and_tmp_464}, or_tmp_1672);
  assign and_4566_cse = and_dcpl_3993 & and_dcpl_4099;
  assign and_4573_cse = (~((~(or_dcpl_857 | or_dcpl_865)) | if_7_equal_svs_st_1))
      & and_dcpl_3998 & and_dcpl_4104;
  assign and_4581_cse = ((else_7_if_1_acc_tmp[2]) | (~ (else_7_if_1_acc_tmp[0]))
      | (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[1]) | (~ else_7_equal_tmp)
      | if_7_equal_tmp) & ((~ (else_7_if_1_div_9cyc[0])) | (else_7_if_1_div_9cyc[1])
      | (else_7_if_1_div_9cyc[3]) | (else_7_if_1_div_9cyc[2]) | (~ else_7_equal_svs_st_1)
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4006 & and_dcpl_4111;
  assign and_4589_cse = or_tmp_1671 & mux_375_cse & and_dcpl_4121 & and_dcpl_4010;
  assign and_4598_cse = or_tmp_1675 & or_tmp_1671 & mux_375_cse & and_dcpl_4020 &
      and_dcpl_4125;
  assign and_4608_cse = or_tmp_1680 & or_tmp_1675 & or_tmp_1671 & mux_375_cse & and_dcpl_4027
      & and_dcpl_868 & (else_7_if_1_div_9cyc_st_5[0]);
  assign and_4619_cse = or_tmp_1686 & or_tmp_1680 & or_tmp_1675 & or_tmp_1671 & mux_375_cse
      & and_dcpl_4034 & and_dcpl_4139;
  assign and_4631_cse = or_tmp_1693 & or_tmp_1686 & or_tmp_1680 & or_tmp_1675 & mux_379_cse
      & and_dcpl_4041 & and_dcpl_4146;
  assign and_4637_cse = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (~ (else_7_if_1_div_9cyc_st_7[0])) | (else_7_if_1_div_9cyc_st_7[1]) | (else_7_if_1_div_9cyc_st_7[2])
      | (else_7_if_1_div_9cyc_st_7[3])) & or_tmp_1693 & or_tmp_1686 & or_tmp_1680
      & or_tmp_1675 & mux_379_cse;
  assign div_mgc_div_20_b = {reg_div_mgc_div_20_b_tmp , 16'b0};
  assign div_mgc_div_20_a = {reg_div_mgc_div_20_a_tmp , 32'b0};
  assign mux_387_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_1753)))
      , or_tmp_1753}, or_tmp_1752);
  assign mux_391_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_507)))
      , and_tmp_507}, or_tmp_1752);
  assign and_4717_cse = and_dcpl_4209 & and_dcpl_3991;
  assign and_4724_cse = (~((~(or_dcpl_877 | or_dcpl_855)) | if_7_equal_svs_st_1))
      & and_dcpl_3998 & and_dcpl_4212;
  assign and_4732_cse = ((else_7_if_1_acc_tmp[2]) | (else_7_if_1_acc_tmp[0]) | (else_7_if_1_acc_tmp[3])
      | (~ (else_7_if_1_acc_tmp[1])) | (~ else_7_equal_tmp) | if_7_equal_tmp) & ((else_7_if_1_div_9cyc[0])
      | (~ (else_7_if_1_div_9cyc[1])) | (else_7_if_1_div_9cyc[3]) | (else_7_if_1_div_9cyc[2])
      | (~ else_7_equal_svs_st_1) | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4006
      & and_dcpl_4219;
  assign and_4740_cse = or_tmp_1751 & mux_387_cse & and_dcpl_4013 & and_dcpl_4226;
  assign and_4749_cse = or_tmp_1755 & or_tmp_1751 & mux_387_cse & and_dcpl_4020 &
      and_dcpl_4233;
  assign and_4759_cse = or_tmp_1760 & or_tmp_1755 & or_tmp_1751 & mux_387_cse & and_dcpl_4027
      & and_dcpl_892 & (~ (else_7_if_1_div_9cyc_st_5[0]));
  assign and_4770_cse = or_tmp_1766 & or_tmp_1760 & or_tmp_1755 & or_tmp_1751 & mux_387_cse
      & and_dcpl_4034 & and_dcpl_4247;
  assign and_4782_cse = or_tmp_1773 & or_tmp_1766 & or_tmp_1760 & or_tmp_1755 & mux_391_cse
      & and_dcpl_4041 & and_dcpl_4254;
  assign and_4788_cse = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (else_7_if_1_div_9cyc_st_7[0]) | (~ (else_7_if_1_div_9cyc_st_7[1])) | (else_7_if_1_div_9cyc_st_7[2])
      | (else_7_if_1_div_9cyc_st_7[3])) & or_tmp_1773 & or_tmp_1766 & or_tmp_1760
      & or_tmp_1755 & mux_391_cse;
  assign div_mgc_div_21_b = {reg_div_mgc_div_21_b_tmp , 16'b0};
  assign div_mgc_div_21_a = {reg_div_mgc_div_21_a_tmp , 32'b0};
  assign mux_399_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_1833)))
      , or_tmp_1833}, or_tmp_1832);
  assign mux_403_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_550)))
      , and_tmp_550}, or_tmp_1832);
  assign and_4868_cse = and_dcpl_4209 & and_dcpl_4099;
  assign and_4875_cse = (~((~(or_dcpl_877 | or_dcpl_865)) | if_7_equal_svs_st_1))
      & and_dcpl_3998 & and_dcpl_4320;
  assign and_4883_cse = ((else_7_if_1_acc_tmp[2]) | (~ (else_7_if_1_acc_tmp[0]))
      | (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[1])) | (~ else_7_equal_tmp)
      | if_7_equal_tmp) & ((~ (else_7_if_1_div_9cyc[0])) | (~ (else_7_if_1_div_9cyc[1]))
      | (else_7_if_1_div_9cyc[3]) | (else_7_if_1_div_9cyc[2]) | (~ else_7_equal_svs_st_1)
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4006 & and_dcpl_4327;
  assign and_4891_cse = or_tmp_1831 & mux_399_cse & and_dcpl_4121 & and_dcpl_4226;
  assign and_4900_cse = or_tmp_1835 & or_tmp_1831 & mux_399_cse & and_dcpl_4020 &
      and_dcpl_4341;
  assign and_4910_cse = or_tmp_1840 & or_tmp_1835 & or_tmp_1831 & mux_399_cse & and_dcpl_4027
      & and_dcpl_892 & (else_7_if_1_div_9cyc_st_5[0]);
  assign and_4921_cse = or_tmp_1846 & or_tmp_1840 & or_tmp_1835 & or_tmp_1831 & mux_399_cse
      & and_dcpl_4034 & and_dcpl_4355;
  assign and_4933_cse = or_tmp_1853 & or_tmp_1846 & or_tmp_1840 & or_tmp_1835 & mux_403_cse
      & and_dcpl_4041 & and_dcpl_4362;
  assign and_4939_cse = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (~ (else_7_if_1_div_9cyc_st_7[0])) | (~ (else_7_if_1_div_9cyc_st_7[1])) |
      (else_7_if_1_div_9cyc_st_7[2]) | (else_7_if_1_div_9cyc_st_7[3])) & or_tmp_1853
      & or_tmp_1846 & or_tmp_1840 & or_tmp_1835 & mux_403_cse;
  assign div_mgc_div_22_b = {reg_div_mgc_div_22_b_tmp , 16'b0};
  assign div_mgc_div_22_a = {reg_div_mgc_div_22_a_tmp , 32'b0};
  assign mux_411_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_1913)))
      , or_tmp_1913}, or_tmp_1912);
  assign mux_415_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_593)))
      , and_tmp_593}, or_tmp_1912);
  assign and_5019_cse = and_dcpl_3993 & and_dcpl_4423;
  assign and_5026_cse = (~((~(or_dcpl_857 | or_dcpl_895)) | if_7_equal_svs_st_1))
      & and_dcpl_4430 & and_dcpl_3996;
  assign and_5034_cse = ((~ (else_7_if_1_acc_tmp[2])) | (else_7_if_1_acc_tmp[0])
      | (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[1]) | (~ else_7_equal_tmp)
      | if_7_equal_tmp) & ((else_7_if_1_div_9cyc[0]) | (else_7_if_1_div_9cyc[1])
      | (else_7_if_1_div_9cyc[3]) | (~ (else_7_if_1_div_9cyc[2])) | (~ else_7_equal_svs_st_1)
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4438 & and_dcpl_4003;
  assign and_5042_cse = or_tmp_1911 & mux_411_cse & and_dcpl_4013 & and_dcpl_4442;
  assign and_5051_cse = or_tmp_1915 & or_tmp_1911 & mux_411_cse & and_dcpl_4452 &
      and_dcpl_4017;
  assign and_5061_cse = or_tmp_1920 & or_tmp_1915 & or_tmp_1911 & mux_411_cse & and_dcpl_4027
      & and_dcpl_916 & (~ (else_7_if_1_div_9cyc_st_5[0]));
  assign and_5072_cse = or_tmp_1926 & or_tmp_1920 & or_tmp_1915 & or_tmp_1911 & mux_411_cse
      & and_dcpl_4466 & and_dcpl_4031;
  assign and_5084_cse = or_tmp_1933 & or_tmp_1926 & or_tmp_1920 & or_tmp_1915 & mux_415_cse
      & and_dcpl_4473 & and_dcpl_4038;
  assign and_5090_cse = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (else_7_if_1_div_9cyc_st_7[0]) | (else_7_if_1_div_9cyc_st_7[1]) | (~ (else_7_if_1_div_9cyc_st_7[2]))
      | (else_7_if_1_div_9cyc_st_7[3])) & or_tmp_1933 & or_tmp_1926 & or_tmp_1920
      & or_tmp_1915 & mux_415_cse;
  assign div_mgc_div_23_b = {reg_div_mgc_div_23_b_tmp , 16'b0};
  assign div_mgc_div_23_a = {reg_div_mgc_div_23_a_tmp , 32'b0};
  assign mux_423_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_1993)))
      , or_tmp_1993}, or_tmp_1992);
  assign mux_427_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_636)))
      , and_tmp_636}, or_tmp_1992);
  assign and_5170_cse = and_dcpl_3993 & and_dcpl_4531;
  assign and_5177_cse = (~((~(or_dcpl_857 | or_dcpl_905)) | if_7_equal_svs_st_1))
      & and_dcpl_4430 & and_dcpl_4104;
  assign and_5185_cse = ((~ (else_7_if_1_acc_tmp[2])) | (~ (else_7_if_1_acc_tmp[0]))
      | (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[1]) | (~ else_7_equal_tmp)
      | if_7_equal_tmp) & ((~ (else_7_if_1_div_9cyc[0])) | (else_7_if_1_div_9cyc[1])
      | (else_7_if_1_div_9cyc[3]) | (~ (else_7_if_1_div_9cyc[2])) | (~ else_7_equal_svs_st_1)
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4438 & and_dcpl_4111;
  assign and_5193_cse = or_tmp_1991 & mux_423_cse & and_dcpl_4121 & and_dcpl_4442;
  assign and_5202_cse = or_tmp_1995 & or_tmp_1991 & mux_423_cse & and_dcpl_4452 &
      and_dcpl_4125;
  assign and_5212_cse = or_tmp_2000 & or_tmp_1995 & or_tmp_1991 & mux_423_cse & and_dcpl_4027
      & and_dcpl_916 & (else_7_if_1_div_9cyc_st_5[0]);
  assign and_5223_cse = or_tmp_2006 & or_tmp_2000 & or_tmp_1995 & or_tmp_1991 & mux_423_cse
      & and_dcpl_4466 & and_dcpl_4139;
  assign and_5235_cse = or_tmp_2013 & or_tmp_2006 & or_tmp_2000 & or_tmp_1995 & mux_427_cse
      & and_dcpl_4473 & and_dcpl_4146;
  assign and_5241_cse = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (~ (else_7_if_1_div_9cyc_st_7[0])) | (else_7_if_1_div_9cyc_st_7[1]) | (~
      (else_7_if_1_div_9cyc_st_7[2])) | (else_7_if_1_div_9cyc_st_7[3])) & or_tmp_2013
      & or_tmp_2006 & or_tmp_2000 & or_tmp_1995 & mux_427_cse;
  assign div_mgc_div_24_b = {reg_div_mgc_div_24_b_tmp , 16'b0};
  assign div_mgc_div_24_a = {reg_div_mgc_div_24_a_tmp , 32'b0};
  assign mux_435_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_2073)))
      , or_tmp_2073}, or_tmp_2072);
  assign mux_439_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_679)))
      , and_tmp_679}, or_tmp_2072);
  assign and_5321_cse = and_dcpl_4209 & and_dcpl_4423;
  assign and_5328_cse = (~((~(or_dcpl_877 | or_dcpl_895)) | if_7_equal_svs_st_1))
      & and_dcpl_4430 & and_dcpl_4212;
  assign and_5336_cse = ((~ (else_7_if_1_acc_tmp[2])) | (else_7_if_1_acc_tmp[0])
      | (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[1])) | (~ else_7_equal_tmp)
      | if_7_equal_tmp) & ((else_7_if_1_div_9cyc[0]) | (~ (else_7_if_1_div_9cyc[1]))
      | (else_7_if_1_div_9cyc[3]) | (~ (else_7_if_1_div_9cyc[2])) | (~ else_7_equal_svs_st_1)
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4438 & and_dcpl_4219;
  assign and_5344_cse = or_tmp_2071 & mux_435_cse & and_dcpl_4013 & and_dcpl_4658;
  assign and_5353_cse = or_tmp_2075 & or_tmp_2071 & mux_435_cse & and_dcpl_4452 &
      and_dcpl_4233;
  assign and_5363_cse = or_tmp_2080 & or_tmp_2075 & or_tmp_2071 & mux_435_cse & and_dcpl_4027
      & and_dcpl_940 & (~ (else_7_if_1_div_9cyc_st_5[0]));
  assign and_5374_cse = or_tmp_2086 & or_tmp_2080 & or_tmp_2075 & or_tmp_2071 & mux_435_cse
      & and_dcpl_4466 & and_dcpl_4247;
  assign and_5386_cse = or_tmp_2093 & or_tmp_2086 & or_tmp_2080 & or_tmp_2075 & mux_439_cse
      & and_dcpl_4473 & and_dcpl_4254;
  assign and_5392_cse = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (else_7_if_1_div_9cyc_st_7[0]) | (~ (else_7_if_1_div_9cyc_st_7[1])) | (~
      (else_7_if_1_div_9cyc_st_7[2])) | (else_7_if_1_div_9cyc_st_7[3])) & or_tmp_2093
      & or_tmp_2086 & or_tmp_2080 & or_tmp_2075 & mux_439_cse;
  assign div_mgc_div_25_b = {reg_div_mgc_div_25_b_tmp , 16'b0};
  assign div_mgc_div_25_a = {reg_div_mgc_div_25_a_tmp , 32'b0};
  assign mux_447_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_2153)))
      , or_tmp_2153}, or_tmp_2152);
  assign mux_451_cse = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_722)))
      , and_tmp_722}, or_tmp_2152);
  assign and_5472_cse = and_dcpl_4209 & and_dcpl_4531;
  assign and_5479_cse = (~((~(or_dcpl_877 | or_dcpl_905)) | if_7_equal_svs_st_1))
      & and_dcpl_4430 & and_dcpl_4320;
  assign and_5487_cse = ((~ (else_7_if_1_acc_tmp[2])) | (~ (else_7_if_1_acc_tmp[0]))
      | (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[1])) | (~ else_7_equal_tmp)
      | if_7_equal_tmp) & (~((else_7_if_1_div_9cyc[0]) & (else_7_if_1_div_9cyc[1])
      & (~ (else_7_if_1_div_9cyc[3])) & (else_7_if_1_div_9cyc[2]) & else_7_equal_svs_st_1
      & main_stage_0_2 & (~ if_7_equal_svs_st_1))) & and_dcpl_4438 & and_dcpl_4327;
  assign and_5495_cse = or_tmp_2151 & mux_447_cse & and_dcpl_4121 & and_dcpl_4658;
  assign and_5504_cse = or_tmp_2155 & or_tmp_2151 & mux_447_cse & and_dcpl_4452 &
      and_dcpl_4341;
  assign and_5514_cse = or_tmp_2160 & or_tmp_2155 & or_tmp_2151 & mux_447_cse & and_dcpl_4027
      & and_dcpl_940 & (else_7_if_1_div_9cyc_st_5[0]);
  assign and_5525_cse = or_tmp_2166 & or_tmp_2160 & or_tmp_2155 & or_tmp_2151 & mux_447_cse
      & and_dcpl_4466 & and_dcpl_4355;
  assign and_5537_cse = or_tmp_2173 & or_tmp_2166 & or_tmp_2160 & or_tmp_2155 & mux_451_cse
      & and_dcpl_4473 & and_dcpl_4362;
  assign and_5543_cse = (~(main_stage_0_8 & (~ if_7_equal_svs_st_7) & else_7_equal_svs_st_7
      & (else_7_if_1_div_9cyc_st_7[0]) & (else_7_if_1_div_9cyc_st_7[1]) & (else_7_if_1_div_9cyc_st_7[2])
      & (~ (else_7_if_1_div_9cyc_st_7[3])))) & or_tmp_2173 & or_tmp_2166 & or_tmp_2160
      & or_tmp_2155 & mux_451_cse;
  assign div_mgc_div_26_b = {reg_div_mgc_div_26_b_tmp , 16'b0};
  assign div_mgc_div_26_a = {reg_div_mgc_div_26_a_tmp , 32'b0};
  assign and_5623_cse = and_dcpl_3993 & (else_7_if_1_acc_tmp[3]) & (~ (else_7_if_1_acc_tmp[0]))
      & (~ (else_7_if_1_acc_tmp[2]));
  assign and_5630_cse = (~((~(or_dcpl_857 | or_dcpl_935)) | if_7_equal_svs_st_1))
      & and_dcpl_3998 & (else_7_if_1_div_9cyc[3]) & (~ (else_7_if_1_div_9cyc[1]))
      & (~ (else_7_if_1_div_9cyc[0]));
  assign and_5638_cse = ((else_7_if_1_acc_tmp[2]) | (else_7_if_1_acc_tmp[0]) | (~
      (else_7_if_1_acc_tmp[3])) | (else_7_if_1_acc_tmp[1]) | (~ else_7_equal_tmp)
      | if_7_equal_tmp) & ((else_7_if_1_div_9cyc[0]) | (else_7_if_1_div_9cyc[1])
      | (~ (else_7_if_1_div_9cyc[3])) | (else_7_if_1_div_9cyc[2]) | (~ else_7_equal_svs_st_1)
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4006 & (else_7_if_1_div_9cyc_st_2[3])
      & (~ (else_7_if_1_div_9cyc_st_2[1])) & (~ (else_7_if_1_div_9cyc_st_2[0]));
  assign mux_460_cse = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_2[3]) | (~ mux_tmp_376)))
      , mux_tmp_376}, or_tmp_2231);
  assign and_5645_cse = mux_460_cse & and_dcpl_4013 & (else_7_if_1_div_9cyc_st_3[3])
      & (~ (else_7_if_1_div_9cyc_st_3[1])) & (~ (else_7_if_1_div_9cyc_st_3[2]));
  assign div_mgc_div_b = {reg_div_mgc_div_b_tmp , 16'b0};
  assign div_mgc_div_a = {reg_div_mgc_div_a_tmp , 32'b0};
  assign and_5737_cse = and_dcpl_4966 & and_dcpl_4963;
  assign and_5745_cse = (~((~(or_dcpl_948 | or_dcpl_945)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_4969;
  assign and_5754_cse = ((else_7_else_1_if_acc_tmp[2]) | (else_7_else_1_if_acc_tmp[0])
      | (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[1]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_if_div_9cyc[0]) | (else_7_else_1_if_div_9cyc[2])
      | (else_7_else_1_if_div_9cyc[1]) | (else_7_else_1_if_div_9cyc[3]) | (~ else_7_else_1_equal_svs_1)
      | else_7_equal_svs_st_1 | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4981
      & and_dcpl_2095 & and_dcpl_2094;
  assign mux_509_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_760)))
      , and_tmp_760}, or_tmp_2353);
  assign and_5763_cse = (mux_509_nl) & and_dcpl_4989 & and_dcpl_1723 & and_dcpl_1722;
  assign mux_510_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_762)))
      , and_tmp_762}, or_tmp_2353);
  assign and_5773_cse = (mux_510_nl) & and_dcpl_4997 & and_dcpl_1351 & and_dcpl_1350;
  assign mux_511_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_765)))
      , and_tmp_765}, or_tmp_2353);
  assign and_5784_cse = (mux_511_nl) & and_dcpl_5005 & and_dcpl_979 & and_dcpl_978;
  assign mux_512_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_769)))
      , and_tmp_769}, or_tmp_2353);
  assign and_5796_cse = (mux_512_nl) & and_dcpl_5013 & and_dcpl_607 & and_dcpl_606;
  assign mux_513_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_774)))
      , and_tmp_774}, or_tmp_2353);
  assign and_5809_cse = (mux_513_nl) & and_dcpl_5021 & and_dcpl_235 & and_dcpl_234;
  assign mux_514_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_780)))
      , and_tmp_780}, or_tmp_2353);
  assign div_mgc_div_10_b = {reg_div_mgc_div_10_b_tmp , 16'b0};
  assign div_mgc_div_10_a = {reg_div_mgc_div_10_a_tmp , 32'b0};
  assign and_5904_cse = and_dcpl_4966 & and_dcpl_5087;
  assign and_5912_cse = (~((~(or_dcpl_948 | or_dcpl_957)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_4968 & (else_7_else_1_if_div_9cyc[0]);
  assign and_5921_cse = ((else_7_else_1_if_acc_tmp[2]) | (~ (else_7_else_1_if_acc_tmp[0]))
      | (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[1]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_if_div_9cyc[0]))
      | (else_7_else_1_if_div_9cyc[2]) | (else_7_else_1_if_div_9cyc[1]) | (else_7_else_1_if_div_9cyc[3])
      | (~ else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1 | (~ main_stage_0_2)
      | if_7_equal_svs_st_1) & and_dcpl_4981 & and_dcpl_2095 & and_dcpl_2108;
  assign mux_521_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_803)))
      , and_tmp_803}, or_tmp_2433);
  assign and_5930_cse = (mux_521_nl) & and_dcpl_4989 & and_dcpl_1737 & and_dcpl_1722;
  assign mux_522_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_805)))
      , and_tmp_805}, or_tmp_2433);
  assign and_5940_cse = (mux_522_nl) & and_dcpl_4997 & and_dcpl_1351 & and_dcpl_1364;
  assign mux_523_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_808)))
      , and_tmp_808}, or_tmp_2433);
  assign and_5951_cse = (mux_523_nl) & and_dcpl_5005 & and_dcpl_979 & and_dcpl_992;
  assign mux_524_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_812)))
      , and_tmp_812}, or_tmp_2433);
  assign and_5963_cse = (mux_524_nl) & and_dcpl_5013 & and_dcpl_607 & and_dcpl_620;
  assign mux_525_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_817)))
      , and_tmp_817}, or_tmp_2433);
  assign and_5976_cse = (mux_525_nl) & and_dcpl_5021 & and_dcpl_235 & and_dcpl_248;
  assign mux_526_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_823)))
      , and_tmp_823}, or_tmp_2433);
  assign div_mgc_div_11_b = {reg_div_mgc_div_11_b_tmp , 16'b0};
  assign div_mgc_div_11_a = {reg_div_mgc_div_11_a_tmp , 32'b0};
  assign and_6071_cse = and_dcpl_5214 & and_dcpl_4963;
  assign and_6079_cse = (~((~(or_dcpl_972 | or_dcpl_945)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_5216 & (~ (else_7_else_1_if_div_9cyc[0]));
  assign and_6088_cse = ((else_7_else_1_if_acc_tmp[2]) | (else_7_else_1_if_acc_tmp[0])
      | (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[1])) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_if_div_9cyc[0]) | (else_7_else_1_if_div_9cyc[2])
      | (~ (else_7_else_1_if_div_9cyc[1])) | (else_7_else_1_if_div_9cyc[3]) | (~
      else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1 | (~ main_stage_0_2) | if_7_equal_svs_st_1)
      & and_dcpl_4981 & and_dcpl_2123 & and_dcpl_2094;
  assign mux_533_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_846)))
      , and_tmp_846}, or_tmp_2513);
  assign and_6097_cse = (mux_533_nl) & and_dcpl_4989 & and_dcpl_1723 & and_dcpl_1750;
  assign mux_534_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_848)))
      , and_tmp_848}, or_tmp_2513);
  assign and_6107_cse = (mux_534_nl) & and_dcpl_4997 & and_dcpl_1351 & and_dcpl_1378;
  assign mux_535_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_851)))
      , and_tmp_851}, or_tmp_2513);
  assign and_6118_cse = (mux_535_nl) & and_dcpl_5005 & and_dcpl_979 & and_dcpl_1006;
  assign mux_536_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_855)))
      , and_tmp_855}, or_tmp_2513);
  assign and_6130_cse = (mux_536_nl) & and_dcpl_5013 & and_dcpl_607 & and_dcpl_634;
  assign mux_537_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_860)))
      , and_tmp_860}, or_tmp_2513);
  assign and_6143_cse = (mux_537_nl) & and_dcpl_5021 & and_dcpl_235 & and_dcpl_262;
  assign mux_538_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_866)))
      , and_tmp_866}, or_tmp_2513);
  assign div_mgc_div_12_b = {reg_div_mgc_div_12_b_tmp , 16'b0};
  assign div_mgc_div_12_a = {reg_div_mgc_div_12_a_tmp , 32'b0};
  assign and_6238_cse = and_dcpl_5214 & and_dcpl_5087;
  assign and_6246_cse = (~((~(or_dcpl_972 | or_dcpl_957)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_5216 & (else_7_else_1_if_div_9cyc[0]);
  assign and_6255_cse = ((else_7_else_1_if_acc_tmp[2]) | (~ (else_7_else_1_if_acc_tmp[0]))
      | (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[1])) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_if_div_9cyc[0]))
      | (else_7_else_1_if_div_9cyc[2]) | (~ (else_7_else_1_if_div_9cyc[1])) | (else_7_else_1_if_div_9cyc[3])
      | (~ else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1 | (~ main_stage_0_2)
      | if_7_equal_svs_st_1) & and_dcpl_4981 & and_dcpl_2123 & and_dcpl_2108;
  assign mux_545_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_889)))
      , and_tmp_889}, or_tmp_2593);
  assign and_6264_cse = (mux_545_nl) & and_dcpl_4989 & and_dcpl_1737 & and_dcpl_1750;
  assign mux_546_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_891)))
      , and_tmp_891}, or_tmp_2593);
  assign and_6274_cse = (mux_546_nl) & and_dcpl_4997 & and_dcpl_1351 & and_dcpl_1392;
  assign mux_547_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_894)))
      , and_tmp_894}, or_tmp_2593);
  assign and_6285_cse = (mux_547_nl) & and_dcpl_5005 & and_dcpl_979 & and_dcpl_1020;
  assign mux_548_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_898)))
      , and_tmp_898}, or_tmp_2593);
  assign and_6297_cse = (mux_548_nl) & and_dcpl_5013 & and_dcpl_607 & and_dcpl_648;
  assign mux_549_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_903)))
      , and_tmp_903}, or_tmp_2593);
  assign and_6310_cse = (mux_549_nl) & and_dcpl_5021 & and_dcpl_235 & and_dcpl_276;
  assign mux_550_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_909)))
      , and_tmp_909}, or_tmp_2593);
  assign div_mgc_div_13_b = {reg_div_mgc_div_13_b_tmp , 16'b0};
  assign div_mgc_div_13_a = {reg_div_mgc_div_13_a_tmp , 32'b0};
  assign and_6405_cse = and_dcpl_4966 & and_dcpl_5459;
  assign and_6413_cse = (~((~(or_dcpl_948 | or_dcpl_993)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_5464 & (~ (else_7_else_1_if_div_9cyc[0]));
  assign and_6422_cse = ((~ (else_7_else_1_if_acc_tmp[2])) | (else_7_else_1_if_acc_tmp[0])
      | (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[1]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_if_div_9cyc[0]) | (~
      (else_7_else_1_if_div_9cyc[2])) | (else_7_else_1_if_div_9cyc[1]) | (else_7_else_1_if_div_9cyc[3])
      | (~ else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1 | (~ main_stage_0_2)
      | if_7_equal_svs_st_1) & and_dcpl_4981 & and_dcpl_2095 & and_dcpl_2150;
  assign mux_557_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_932)))
      , and_tmp_932}, or_tmp_2673);
  assign and_6431_cse = (mux_557_nl) & and_dcpl_4989 & and_dcpl_1723 & and_dcpl_1778;
  assign mux_558_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_934)))
      , and_tmp_934}, or_tmp_2673);
  assign and_6441_cse = (mux_558_nl) & and_dcpl_4997 & and_dcpl_1407 & and_dcpl_1350;
  assign mux_559_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_937)))
      , and_tmp_937}, or_tmp_2673);
  assign and_6452_cse = (mux_559_nl) & and_dcpl_5005 & and_dcpl_1035 & and_dcpl_978;
  assign mux_560_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_941)))
      , and_tmp_941}, or_tmp_2673);
  assign and_6464_cse = (mux_560_nl) & and_dcpl_5013 & and_dcpl_663 & and_dcpl_606;
  assign mux_561_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_946)))
      , and_tmp_946}, or_tmp_2673);
  assign and_6477_cse = (mux_561_nl) & and_dcpl_5021 & and_dcpl_291 & and_dcpl_234;
  assign mux_562_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_952)))
      , and_tmp_952}, or_tmp_2673);
  assign div_mgc_div_14_b = {reg_div_mgc_div_14_b_tmp , 16'b0};
  assign div_mgc_div_14_a = {reg_div_mgc_div_14_a_tmp , 32'b0};
  assign and_6572_cse = and_dcpl_4966 & and_dcpl_5583;
  assign and_6580_cse = (~((~(or_dcpl_948 | or_dcpl_1005)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_5464 & (else_7_else_1_if_div_9cyc[0]);
  assign and_6589_cse = ((~ (else_7_else_1_if_acc_tmp[2])) | (~ (else_7_else_1_if_acc_tmp[0]))
      | (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[1]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_if_div_9cyc[0]))
      | (~ (else_7_else_1_if_div_9cyc[2])) | (else_7_else_1_if_div_9cyc[1]) | (else_7_else_1_if_div_9cyc[3])
      | (~ else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1 | (~ main_stage_0_2)
      | if_7_equal_svs_st_1) & and_dcpl_4981 & and_dcpl_2095 & and_dcpl_2164;
  assign mux_569_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_975)))
      , and_tmp_975}, or_tmp_2753);
  assign and_6598_cse = (mux_569_nl) & and_dcpl_4989 & and_dcpl_1737 & and_dcpl_1778;
  assign mux_570_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_977)))
      , and_tmp_977}, or_tmp_2753);
  assign and_6608_cse = (mux_570_nl) & and_dcpl_4997 & and_dcpl_1407 & and_dcpl_1364;
  assign mux_571_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_980)))
      , and_tmp_980}, or_tmp_2753);
  assign and_6619_cse = (mux_571_nl) & and_dcpl_5005 & and_dcpl_1035 & and_dcpl_992;
  assign mux_572_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_984)))
      , and_tmp_984}, or_tmp_2753);
  assign and_6631_cse = (mux_572_nl) & and_dcpl_5013 & and_dcpl_663 & and_dcpl_620;
  assign mux_573_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_989)))
      , and_tmp_989}, or_tmp_2753);
  assign and_6644_cse = (mux_573_nl) & and_dcpl_5021 & and_dcpl_291 & and_dcpl_248;
  assign mux_574_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_995)))
      , and_tmp_995}, or_tmp_2753);
  assign div_mgc_div_15_b = {reg_div_mgc_div_15_b_tmp , 16'b0};
  assign div_mgc_div_15_a = {reg_div_mgc_div_15_a_tmp , 32'b0};
  assign and_6739_cse = and_dcpl_5214 & and_dcpl_5459;
  assign and_6747_cse = (~((~(or_dcpl_972 | or_dcpl_993)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_5712 & (~ (else_7_else_1_if_div_9cyc[0]));
  assign and_6756_cse = ((~ (else_7_else_1_if_acc_tmp[2])) | (else_7_else_1_if_acc_tmp[0])
      | (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[1])) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_if_div_9cyc[0]) | (~
      (else_7_else_1_if_div_9cyc[2])) | (~ (else_7_else_1_if_div_9cyc[1])) | (else_7_else_1_if_div_9cyc[3])
      | (~ else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1 | (~ main_stage_0_2)
      | if_7_equal_svs_st_1) & and_dcpl_4981 & and_dcpl_2123 & and_dcpl_2150;
  assign mux_581_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1018)))
      , and_tmp_1018}, or_tmp_2833);
  assign and_6765_cse = (mux_581_nl) & and_dcpl_4989 & and_dcpl_1723 & and_dcpl_1806;
  assign mux_582_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1020)))
      , and_tmp_1020}, or_tmp_2833);
  assign and_6775_cse = (mux_582_nl) & and_dcpl_4997 & and_dcpl_1407 & and_dcpl_1378;
  assign mux_583_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1023)))
      , and_tmp_1023}, or_tmp_2833);
  assign and_6786_cse = (mux_583_nl) & and_dcpl_5005 & and_dcpl_1035 & and_dcpl_1006;
  assign mux_584_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1027)))
      , and_tmp_1027}, or_tmp_2833);
  assign and_6798_cse = (mux_584_nl) & and_dcpl_5013 & and_dcpl_663 & and_dcpl_634;
  assign mux_585_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1032)))
      , and_tmp_1032}, or_tmp_2833);
  assign and_6811_cse = (mux_585_nl) & and_dcpl_5021 & and_dcpl_291 & and_dcpl_262;
  assign mux_586_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1038)))
      , and_tmp_1038}, or_tmp_2833);
  assign div_mgc_div_16_b = {reg_div_mgc_div_16_b_tmp , 16'b0};
  assign div_mgc_div_16_a = {reg_div_mgc_div_16_a_tmp , 32'b0};
  assign and_6906_cse = and_dcpl_5214 & and_dcpl_5583;
  assign and_6914_cse = (~((~(or_dcpl_972 | or_dcpl_1005)) | if_7_equal_svs_st_1))
      & and_dcpl_4972 & and_dcpl_5712 & (else_7_else_1_if_div_9cyc[0]);
  assign and_6923_cse = ((~ (else_7_else_1_if_acc_tmp[2])) | (~ (else_7_else_1_if_acc_tmp[0]))
      | (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[1])) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_if_div_9cyc[0]))
      | (~ (else_7_else_1_if_div_9cyc[2])) | (~ (else_7_else_1_if_div_9cyc[1])) |
      (else_7_else_1_if_div_9cyc[3]) | (~ else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_dcpl_4981 & and_dcpl_2123
      & and_dcpl_2164;
  assign mux_593_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1061)))
      , and_tmp_1061}, or_tmp_2913);
  assign and_6932_cse = (mux_593_nl) & and_dcpl_4989 & and_dcpl_1737 & and_dcpl_1806;
  assign mux_594_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1063)))
      , and_tmp_1063}, or_tmp_2913);
  assign and_6942_cse = (mux_594_nl) & and_dcpl_4997 & and_dcpl_1407 & and_dcpl_1392;
  assign mux_595_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1066)))
      , and_tmp_1066}, or_tmp_2913);
  assign and_6953_cse = (mux_595_nl) & and_dcpl_5005 & and_dcpl_1035 & and_dcpl_1020;
  assign mux_596_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1070)))
      , and_tmp_1070}, or_tmp_2913);
  assign and_6965_cse = (mux_596_nl) & and_dcpl_5013 & and_dcpl_663 & and_dcpl_648;
  assign mux_597_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1075)))
      , and_tmp_1075}, or_tmp_2913);
  assign and_6978_cse = (mux_597_nl) & and_dcpl_5021 & and_dcpl_291 & and_dcpl_276;
  assign mux_598_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1081)))
      , and_tmp_1081}, or_tmp_2913);
  assign div_mgc_div_17_b = {reg_div_mgc_div_17_b_tmp , 16'b0};
  assign div_mgc_div_17_a = {reg_div_mgc_div_17_a_tmp , 32'b0};
  assign and_7073_cse = and_dcpl_4966 & (else_7_else_1_if_acc_tmp[3]) & (~ (else_7_else_1_if_acc_tmp[0]))
      & (~ (else_7_else_1_if_acc_tmp[2]));
  assign and_7081_cse = (~((~(or_dcpl_948 | or_dcpl_1041)) | if_7_equal_svs_st_1))
      & and_dcpl_4971 & else_7_else_1_equal_svs_1 & (else_7_else_1_if_div_9cyc[3])
      & and_dcpl_4969;
  assign and_7090_cse = ((else_7_else_1_if_acc_tmp[2]) | (else_7_else_1_if_acc_tmp[0])
      | (~ (else_7_else_1_if_acc_tmp[3])) | (else_7_else_1_if_acc_tmp[1]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_if_div_9cyc[0]) | (else_7_else_1_if_div_9cyc[2])
      | (else_7_else_1_if_div_9cyc[1]) | (~ (else_7_else_1_if_div_9cyc[3])) | (~
      else_7_else_1_equal_svs_1) | else_7_equal_svs_st_1 | (~ main_stage_0_2) | if_7_equal_svs_st_1)
      & and_dcpl_4981 & (else_7_else_1_if_div_9cyc_st_2[3]) & (~ (else_7_else_1_if_div_9cyc_st_2[1]))
      & and_dcpl_2094;
  assign mux_605_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ and_tmp_1104)))
      , and_tmp_1104}, or_tmp_2993);
  assign and_7099_cse = (mux_605_nl) & and_dcpl_4989 & (~ (else_7_else_1_if_div_9cyc_st_3[0]))
      & (else_7_else_1_if_div_9cyc_st_3[3]) & and_dcpl_1722;
  assign div_mgc_div_18_b = {reg_div_mgc_div_18_b_tmp , 16'b0};
  assign div_mgc_div_18_a = {reg_div_mgc_div_18_a_tmp , 32'b0};
  assign and_7204_cse = and_dcpl_6082 & and_dcpl_6079;
  assign and_7212_cse = (~((~(or_dcpl_1056 | or_dcpl_1053)) | if_7_equal_svs_st_1))
      & and_dcpl_6088 & and_dcpl_6085;
  assign and_7221_cse = ((else_7_else_1_else_acc_tmp[2]) | (else_7_else_1_else_acc_tmp[0])
      | (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[1]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_else_div_9cyc[0]) |
      (else_7_else_1_else_div_9cyc[1]) | (else_7_else_1_else_div_9cyc[3]) | (else_7_else_1_else_div_9cyc[2])
      | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1 | (~ main_stage_0_2) |
      if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2224 & and_dcpl_2223;
  assign and_7231_cse = or_tmp_3115 & or_tmp_3116 & or_tmp_3117 & and_1990_cse &
      and_dcpl_1852 & and_dcpl_1851;
  assign and_7242_cse = or_tmp_3115 & or_tmp_3117 & or_tmp_3116 & or_tmp_3121 & and_1618_cse
      & and_dcpl_1480 & and_dcpl_1479;
  assign and_7254_cse = or_tmp_3115 & or_tmp_3123 & or_tmp_3121 & and_tmp_1116 &
      and_1246_cse & and_dcpl_1108 & and_dcpl_1107;
  assign and_7267_cse = or_tmp_3115 & or_tmp_3128 & or_tmp_3123 & or_tmp_3121 & and_tmp_1116
      & and_874_cse & and_dcpl_736 & and_dcpl_735;
  assign and_7281_cse = or_tmp_3115 & or_tmp_3134 & or_tmp_3128 & or_tmp_3123 & or_tmp_3121
      & and_tmp_1116 & and_502_cse & and_dcpl_364 & and_dcpl_363;
  assign and_7288_cse = or_tmp_3115 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (else_7_else_1_else_div_9cyc_st_7[0])
      | (else_7_else_1_else_div_9cyc_st_7[1]) | (else_7_else_1_else_div_9cyc_st_7[2])
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3116 & or_tmp_3134 & or_tmp_3128
      & or_tmp_3123 & or_tmp_3121 & or_tmp_3117;
  assign div_mgc_div_1_b = {reg_div_mgc_div_1_b_tmp , 16'b0};
  assign div_mgc_div_1_a = {reg_div_mgc_div_1_a_tmp , 32'b0};
  assign and_7383_cse = and_dcpl_6082 & and_dcpl_6203;
  assign and_7391_cse = (~((~(or_dcpl_1056 | or_dcpl_1065)) | if_7_equal_svs_st_1))
      & and_dcpl_6088 & and_dcpl_6209;
  assign and_7400_cse = ((else_7_else_1_else_acc_tmp[2]) | (~ (else_7_else_1_else_acc_tmp[0]))
      | (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[1]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_else_div_9cyc[0]))
      | (else_7_else_1_else_div_9cyc[1]) | (else_7_else_1_else_div_9cyc[3]) | (else_7_else_1_else_div_9cyc[2])
      | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1 | (~ main_stage_0_2) |
      if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2224 & and_dcpl_2237;
  assign and_7410_cse = or_tmp_3183 & or_tmp_3184 & or_tmp_3185 & and_1990_cse &
      and_dcpl_1852 & and_dcpl_1865;
  assign and_7421_cse = or_tmp_3183 & or_tmp_3185 & or_tmp_3184 & or_tmp_3189 & and_1618_cse
      & and_dcpl_1480 & and_dcpl_1493;
  assign and_7433_cse = or_tmp_3183 & or_tmp_3191 & or_tmp_3189 & and_tmp_1171 &
      and_1246_cse & and_dcpl_1108 & and_dcpl_1121;
  assign and_7446_cse = or_tmp_3183 & or_tmp_3196 & or_tmp_3191 & or_tmp_3189 & and_tmp_1171
      & and_874_cse & and_dcpl_736 & and_dcpl_749;
  assign and_7460_cse = or_tmp_3183 & or_tmp_3202 & or_tmp_3196 & or_tmp_3191 & or_tmp_3189
      & and_tmp_1171 & and_502_cse & and_dcpl_364 & and_dcpl_377;
  assign and_7467_cse = or_tmp_3183 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (~ (else_7_else_1_else_div_9cyc_st_7[0]))
      | (else_7_else_1_else_div_9cyc_st_7[1]) | (else_7_else_1_else_div_9cyc_st_7[2])
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3184 & or_tmp_3202 & or_tmp_3196
      & or_tmp_3191 & or_tmp_3189 & or_tmp_3185;
  assign div_mgc_div_2_b = {reg_div_mgc_div_2_b_tmp , 16'b0};
  assign div_mgc_div_2_a = {reg_div_mgc_div_2_a_tmp , 32'b0};
  assign and_7562_cse = and_dcpl_6330 & and_dcpl_6079;
  assign and_7570_cse = (~((~(or_dcpl_1080 | or_dcpl_1053)) | if_7_equal_svs_st_1))
      & and_dcpl_6088 & and_dcpl_6333;
  assign and_7579_cse = ((else_7_else_1_else_acc_tmp[2]) | (else_7_else_1_else_acc_tmp[0])
      | (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[1])) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_else_div_9cyc[0]) |
      (~ (else_7_else_1_else_div_9cyc[1])) | (else_7_else_1_else_div_9cyc[3]) | (else_7_else_1_else_div_9cyc[2])
      | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1 | (~ main_stage_0_2) |
      if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2224 & and_dcpl_2251;
  assign and_7589_cse = or_tmp_3251 & or_tmp_3252 & or_tmp_3253 & and_1990_cse &
      and_dcpl_1852 & and_dcpl_1879;
  assign and_7600_cse = or_tmp_3251 & or_tmp_3253 & or_tmp_3252 & or_tmp_3257 & and_1618_cse
      & and_dcpl_1480 & and_dcpl_1507;
  assign and_7612_cse = or_tmp_3251 & or_tmp_3259 & or_tmp_3257 & and_tmp_1226 &
      and_1246_cse & and_dcpl_1108 & and_dcpl_1135;
  assign and_7625_cse = or_tmp_3251 & or_tmp_3264 & or_tmp_3259 & or_tmp_3257 & and_tmp_1226
      & and_874_cse & and_dcpl_736 & and_dcpl_763;
  assign and_7639_cse = or_tmp_3251 & or_tmp_3270 & or_tmp_3264 & or_tmp_3259 & or_tmp_3257
      & and_tmp_1226 & and_502_cse & and_dcpl_364 & and_dcpl_391;
  assign and_7646_cse = or_tmp_3251 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (else_7_else_1_else_div_9cyc_st_7[0])
      | (~ (else_7_else_1_else_div_9cyc_st_7[1])) | (else_7_else_1_else_div_9cyc_st_7[2])
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3252 & or_tmp_3270 & or_tmp_3264
      & or_tmp_3259 & or_tmp_3257 & or_tmp_3253;
  assign div_mgc_div_3_b = {reg_div_mgc_div_3_b_tmp , 16'b0};
  assign div_mgc_div_3_a = {reg_div_mgc_div_3_a_tmp , 32'b0};
  assign and_7741_cse = and_dcpl_6330 & and_dcpl_6203;
  assign and_7749_cse = (~((~(or_dcpl_1080 | or_dcpl_1065)) | if_7_equal_svs_st_1))
      & and_dcpl_6088 & and_dcpl_6457;
  assign and_7758_cse = ((else_7_else_1_else_acc_tmp[2]) | (~ (else_7_else_1_else_acc_tmp[0]))
      | (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[1])) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_else_div_9cyc[0]))
      | (~ (else_7_else_1_else_div_9cyc[1])) | (else_7_else_1_else_div_9cyc[3]) |
      (else_7_else_1_else_div_9cyc[2]) | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2224
      & and_dcpl_2265;
  assign and_7768_cse = or_tmp_3319 & or_tmp_3320 & or_tmp_3321 & and_1990_cse &
      and_dcpl_1852 & and_dcpl_1893;
  assign and_7779_cse = or_tmp_3319 & or_tmp_3321 & or_tmp_3320 & or_tmp_3325 & and_1618_cse
      & and_dcpl_1480 & and_dcpl_1521;
  assign and_7791_cse = or_tmp_3319 & or_tmp_3327 & or_tmp_3325 & and_tmp_1281 &
      and_1246_cse & and_dcpl_1108 & and_dcpl_1149;
  assign and_7804_cse = or_tmp_3319 & or_tmp_3332 & or_tmp_3327 & or_tmp_3325 & and_tmp_1281
      & and_874_cse & and_dcpl_736 & and_dcpl_777;
  assign and_7818_cse = or_tmp_3319 & or_tmp_3338 & or_tmp_3332 & or_tmp_3327 & or_tmp_3325
      & and_tmp_1281 & and_502_cse & and_dcpl_364 & and_dcpl_405;
  assign and_7825_cse = or_tmp_3319 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (~ (else_7_else_1_else_div_9cyc_st_7[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_7[1])) | (else_7_else_1_else_div_9cyc_st_7[2])
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3320 & or_tmp_3338 & or_tmp_3332
      & or_tmp_3327 & or_tmp_3325 & or_tmp_3321;
  assign div_mgc_div_4_b = {reg_div_mgc_div_4_b_tmp , 16'b0};
  assign div_mgc_div_4_a = {reg_div_mgc_div_4_a_tmp , 32'b0};
  assign and_7920_cse = and_dcpl_6082 & and_dcpl_6575;
  assign and_7928_cse = (~((~(or_dcpl_1056 | or_dcpl_1101)) | if_7_equal_svs_st_1))
      & and_dcpl_6584 & and_dcpl_6085;
  assign and_7937_cse = ((~ (else_7_else_1_else_acc_tmp[2])) | (else_7_else_1_else_acc_tmp[0])
      | (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[1]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_else_div_9cyc[0]) |
      (else_7_else_1_else_div_9cyc[1]) | (else_7_else_1_else_div_9cyc[3]) | (~ (else_7_else_1_else_div_9cyc[2]))
      | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1 | (~ main_stage_0_2) |
      if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2280 & and_dcpl_2223;
  assign and_7947_cse = or_tmp_3387 & or_tmp_3388 & or_tmp_3389 & and_1990_cse &
      and_dcpl_1908 & and_dcpl_1851;
  assign and_7958_cse = or_tmp_3387 & or_tmp_3389 & or_tmp_3388 & or_tmp_3393 & and_1618_cse
      & and_dcpl_1536 & and_dcpl_1479;
  assign and_7970_cse = or_tmp_3387 & or_tmp_3395 & or_tmp_3393 & and_tmp_1336 &
      and_1246_cse & and_dcpl_1164 & and_dcpl_1107;
  assign and_7983_cse = or_tmp_3387 & or_tmp_3400 & or_tmp_3395 & or_tmp_3393 & and_tmp_1336
      & and_874_cse & and_dcpl_792 & and_dcpl_735;
  assign and_7997_cse = or_tmp_3387 & or_tmp_3406 & or_tmp_3400 & or_tmp_3395 & or_tmp_3393
      & and_tmp_1336 & and_502_cse & and_dcpl_420 & and_dcpl_363;
  assign and_8004_cse = or_tmp_3387 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (else_7_else_1_else_div_9cyc_st_7[0])
      | (else_7_else_1_else_div_9cyc_st_7[1]) | (~ (else_7_else_1_else_div_9cyc_st_7[2]))
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3388 & or_tmp_3406 & or_tmp_3400
      & or_tmp_3395 & or_tmp_3393 & or_tmp_3389;
  assign div_mgc_div_5_b = {reg_div_mgc_div_5_b_tmp , 16'b0};
  assign div_mgc_div_5_a = {reg_div_mgc_div_5_a_tmp , 32'b0};
  assign and_8099_cse = and_dcpl_6082 & and_dcpl_6699;
  assign and_8107_cse = (~((~(or_dcpl_1056 | or_dcpl_1113)) | if_7_equal_svs_st_1))
      & and_dcpl_6584 & and_dcpl_6209;
  assign and_8116_cse = ((~ (else_7_else_1_else_acc_tmp[2])) | (~ (else_7_else_1_else_acc_tmp[0]))
      | (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[1]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_else_div_9cyc[0]))
      | (else_7_else_1_else_div_9cyc[1]) | (else_7_else_1_else_div_9cyc[3]) | (~
      (else_7_else_1_else_div_9cyc[2])) | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2280
      & and_dcpl_2237;
  assign and_8126_cse = or_tmp_3455 & or_tmp_3456 & or_tmp_3457 & and_1990_cse &
      and_dcpl_1908 & and_dcpl_1865;
  assign and_8137_cse = or_tmp_3455 & or_tmp_3457 & or_tmp_3456 & or_tmp_3461 & and_1618_cse
      & and_dcpl_1536 & and_dcpl_1493;
  assign and_8149_cse = or_tmp_3455 & or_tmp_3463 & or_tmp_3461 & and_tmp_1391 &
      and_1246_cse & and_dcpl_1164 & and_dcpl_1121;
  assign and_8162_cse = or_tmp_3455 & or_tmp_3468 & or_tmp_3463 & or_tmp_3461 & and_tmp_1391
      & and_874_cse & and_dcpl_792 & and_dcpl_749;
  assign and_8176_cse = or_tmp_3455 & or_tmp_3474 & or_tmp_3468 & or_tmp_3463 & or_tmp_3461
      & and_tmp_1391 & and_502_cse & and_dcpl_420 & and_dcpl_377;
  assign and_8183_cse = or_tmp_3455 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (~ (else_7_else_1_else_div_9cyc_st_7[0]))
      | (else_7_else_1_else_div_9cyc_st_7[1]) | (~ (else_7_else_1_else_div_9cyc_st_7[2]))
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3456 & or_tmp_3474 & or_tmp_3468
      & or_tmp_3463 & or_tmp_3461 & or_tmp_3457;
  assign div_mgc_div_6_b = {reg_div_mgc_div_6_b_tmp , 16'b0};
  assign div_mgc_div_6_a = {reg_div_mgc_div_6_a_tmp , 32'b0};
  assign and_8278_cse = and_dcpl_6330 & and_dcpl_6575;
  assign and_8286_cse = (~((~(or_dcpl_1080 | or_dcpl_1101)) | if_7_equal_svs_st_1))
      & and_dcpl_6584 & and_dcpl_6333;
  assign and_8295_cse = ((~ (else_7_else_1_else_acc_tmp[2])) | (else_7_else_1_else_acc_tmp[0])
      | (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[1])) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_else_div_9cyc[0]) |
      (~ (else_7_else_1_else_div_9cyc[1])) | (else_7_else_1_else_div_9cyc[3]) | (~
      (else_7_else_1_else_div_9cyc[2])) | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2280
      & and_dcpl_2251;
  assign and_8305_cse = or_tmp_3523 & or_tmp_3524 & or_tmp_3525 & and_1990_cse &
      and_dcpl_1908 & and_dcpl_1879;
  assign and_8316_cse = or_tmp_3523 & or_tmp_3525 & or_tmp_3524 & or_tmp_3529 & and_1618_cse
      & and_dcpl_1536 & and_dcpl_1507;
  assign and_8328_cse = or_tmp_3523 & or_tmp_3531 & or_tmp_3529 & and_tmp_1446 &
      and_1246_cse & and_dcpl_1164 & and_dcpl_1135;
  assign and_8341_cse = or_tmp_3523 & or_tmp_3536 & or_tmp_3531 & or_tmp_3529 & and_tmp_1446
      & and_874_cse & and_dcpl_792 & and_dcpl_763;
  assign and_8355_cse = or_tmp_3523 & or_tmp_3542 & or_tmp_3536 & or_tmp_3531 & or_tmp_3529
      & and_tmp_1446 & and_502_cse & and_dcpl_420 & and_dcpl_391;
  assign and_8362_cse = or_tmp_3523 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (else_7_else_1_else_div_9cyc_st_7[0])
      | (~ (else_7_else_1_else_div_9cyc_st_7[1])) | (~ (else_7_else_1_else_div_9cyc_st_7[2]))
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3524 & or_tmp_3542 & or_tmp_3536
      & or_tmp_3531 & or_tmp_3529 & or_tmp_3525;
  assign div_mgc_div_7_b = {reg_div_mgc_div_7_b_tmp , 16'b0};
  assign div_mgc_div_7_a = {reg_div_mgc_div_7_a_tmp , 32'b0};
  assign and_8457_cse = and_dcpl_6330 & and_dcpl_6699;
  assign and_8465_cse = (~((~(or_dcpl_1080 | or_dcpl_1113)) | if_7_equal_svs_st_1))
      & and_dcpl_6584 & and_dcpl_6457;
  assign and_8474_cse = ((~ (else_7_else_1_else_acc_tmp[2])) | (~ (else_7_else_1_else_acc_tmp[0]))
      | (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[1])) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((~ (else_7_else_1_else_div_9cyc[0]))
      | (~ (else_7_else_1_else_div_9cyc[1])) | (else_7_else_1_else_div_9cyc[3]) |
      (~ (else_7_else_1_else_div_9cyc[2])) | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1
      | (~ main_stage_0_2) | if_7_equal_svs_st_1) & and_2362_cse & and_dcpl_2280
      & and_dcpl_2265;
  assign and_8484_cse = or_tmp_3591 & or_tmp_3592 & or_tmp_3593 & and_1990_cse &
      and_dcpl_1908 & and_dcpl_1893;
  assign and_8495_cse = or_tmp_3591 & or_tmp_3593 & or_tmp_3592 & or_tmp_3597 & and_1618_cse
      & and_dcpl_1536 & and_dcpl_1521;
  assign and_8507_cse = or_tmp_3591 & or_tmp_3599 & or_tmp_3597 & and_tmp_1501 &
      and_1246_cse & and_dcpl_1164 & and_dcpl_1149;
  assign and_8520_cse = or_tmp_3591 & or_tmp_3604 & or_tmp_3599 & or_tmp_3597 & and_tmp_1501
      & and_874_cse & and_dcpl_792 & and_dcpl_777;
  assign and_8534_cse = or_tmp_3591 & or_tmp_3610 & or_tmp_3604 & or_tmp_3599 & or_tmp_3597
      & and_tmp_1501 & and_502_cse & and_dcpl_420 & and_dcpl_405;
  assign and_8541_cse = or_tmp_3591 & ((~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (~ (else_7_else_1_else_div_9cyc_st_7[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_7[1])) | (~ (else_7_else_1_else_div_9cyc_st_7[2]))
      | (else_7_else_1_else_div_9cyc_st_7[3])) & or_tmp_3592 & or_tmp_3610 & or_tmp_3604
      & or_tmp_3599 & or_tmp_3597 & or_tmp_3593;
  assign div_mgc_div_8_b = {reg_div_mgc_div_8_b_tmp , 16'b0};
  assign div_mgc_div_8_a = {reg_div_mgc_div_8_a_tmp , 32'b0};
  assign and_8636_cse = and_dcpl_6082 & (else_7_else_1_else_acc_tmp[3]) & (~ (else_7_else_1_else_acc_tmp[0]))
      & (~ (else_7_else_1_else_acc_tmp[2]));
  assign and_8644_cse = (~((~(or_dcpl_1056 | or_dcpl_1149)) | if_7_equal_svs_st_1))
      & and_dcpl_6088 & (else_7_else_1_else_div_9cyc[3]) & (~ (else_7_else_1_else_div_9cyc[1]))
      & (~ (else_7_else_1_else_div_9cyc[0]));
  assign and_8653_cse = ((else_7_else_1_else_acc_tmp[2]) | (else_7_else_1_else_acc_tmp[0])
      | (~ (else_7_else_1_else_acc_tmp[3])) | (else_7_else_1_else_acc_tmp[1]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp) & ((else_7_else_1_else_div_9cyc[0]) |
      (else_7_else_1_else_div_9cyc[1]) | (~ (else_7_else_1_else_div_9cyc[3])) | (else_7_else_1_else_div_9cyc[2])
      | else_7_else_1_equal_svs_1 | else_7_equal_svs_st_1 | (~ main_stage_0_2) |
      if_7_equal_svs_st_1) & and_2362_cse & (~ (else_7_else_1_else_div_9cyc_st_2[2]))
      & (else_7_else_1_else_div_9cyc_st_2[3]) & and_dcpl_2223;
  assign and_8663_cse = or_tmp_3659 & or_tmp_3660 & or_tmp_3662 & and_1990_cse &
      (~ (else_7_else_1_else_div_9cyc_st_3[2])) & (else_7_else_1_else_div_9cyc_st_3[3])
      & and_dcpl_1851;
  assign mux_653_nl = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_2[3]) | (~
      and_tmp_1553))) , and_tmp_1553}, or_tmp_3661);
  assign and_8673_cse = or_tmp_3659 & (mux_653_nl) & and_1618_cse & (~ (else_7_else_1_else_div_9cyc_st_4[2]))
      & (else_7_else_1_else_div_9cyc_st_4[3]) & and_dcpl_1479;
  assign div_mgc_div_9_b = {reg_div_mgc_div_9_b_tmp , 16'b0};
  assign div_mgc_div_9_a = {reg_div_mgc_div_9_a_tmp , 32'b0};
  assign and_502_cse = and_dcpl_17 & (~(else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7));
  assign and_874_cse = and_506_cse & (~(else_7_equal_svs_st_6 | else_7_else_1_equal_svs_st_6));
  assign and_1246_cse = and_878_cse & (~(else_7_equal_svs_st_5 | else_7_else_1_equal_svs_st_5));
  assign and_1618_cse = and_1250_cse & (~(else_7_equal_svs_st_4 | else_7_else_1_equal_svs_st_4));
  assign and_1990_cse = and_1622_cse & (~(else_7_equal_svs_st_3 | else_7_else_1_equal_svs_st_3));
  assign and_2362_cse = and_1994_cse & (~(else_7_equal_svs_st_2 | else_7_else_1_equal_svs_st_2));
  assign or_4933_cse = and_9058_cse | or_dcpl_1162 | or_dcpl_1160;
  assign or_4943_cse = and_9058_cse | or_dcpl_1162 | or_dcpl_1170;
  assign or_4953_cse = and_9058_cse | or_dcpl_1162 | or_dcpl_1180;
  assign or_4963_cse = and_9058_cse | or_dcpl_1162 | or_dcpl_1190;
  assign or_4973_cse = and_9058_cse | or_dcpl_1202 | or_dcpl_1160;
  assign or_4983_cse = and_9058_cse | or_dcpl_1202 | or_dcpl_1170;
  assign or_4993_cse = and_9058_cse | or_dcpl_1202 | or_dcpl_1180;
  assign or_5003_cse = and_9058_cse | or_dcpl_1202 | or_dcpl_1190;
  assign or_5013_cse = and_9058_cse | if_7_equal_tmp | (~ (else_7_if_acc_tmp[3]))
      | (else_7_if_acc_tmp[2]) | or_dcpl_1160;
  assign and_9058_cse = (~((mux1h_81_tmp[0]) | (mux1h_81_tmp[1]))) & (~((mux1h_81_tmp[2])
      | (mux1h_81_tmp[3]))) & (~((mux1h_81_tmp[4]) | (mux1h_81_tmp[5]))) & (~((mux1h_81_tmp[6])
      | (mux1h_81_tmp[7]))) & (~((mux1h_81_tmp[8]) | (mux1h_81_tmp[9]))) & (~((mux1h_81_tmp[10])
      | (mux1h_81_tmp[11]))) & (~((mux1h_81_tmp[12]) | (mux1h_81_tmp[13]))) & (~((mux1h_81_tmp[14])
      | (mux1h_81_tmp[15])));
  assign or_5270_cse = or_dcpl_1056 | or_dcpl_1101;
  assign or_5282_cse = or_dcpl_1056 | or_dcpl_1113;
  assign or_5294_cse = or_dcpl_1080 | or_dcpl_1101;
  assign or_5306_cse = or_dcpl_1080 | or_dcpl_1113;
  assign or_5318_cse = or_dcpl_1056 | or_dcpl_1149;
  assign or_5325_cse = and_9058_cse | if_7_equal_tmp;
  assign else_7_acc_2_psp_sg1_sva_1 = MUX_v_16_2_2({(else_7_acc_2_itm[29:14]) , else_7_acc_2_psp_sg1_sva},
      if_7_equal_svs_9);
  assign nl_else_7_acc_2_itm = ({(~ h_2_lpi_dfm_1_sg2_1) , (~ h_2_lpi_dfm_1_sg1_1)
      , (~ h_2_lpi_dfm_4)}) + ({(h_2_lpi_dfm_1_sg2_1[7:0]) , h_2_lpi_dfm_1_sg1_1
      , h_2_lpi_dfm_4 , 4'b1});
  assign else_7_acc_2_itm = nl_else_7_acc_2_itm[29:0];
  assign h_2_sva_duc_mx0 = MUX1HOT_v_30_10_2({(div_mgc_div_19_z[29:0]) , (div_mgc_div_20_z[29:0])
      , (div_mgc_div_21_z[29:0]) , (div_mgc_div_22_z[29:0]) , (div_mgc_div_23_z[29:0])
      , (div_mgc_div_24_z[29:0]) , (div_mgc_div_25_z[29:0]) , (div_mgc_div_26_z[29:0])
      , (div_mgc_div_z[29:0]) , h_2_sva_duc}, {(and_dcpl_2832 & and_dcpl_2831) ,
      (and_dcpl_2835 & and_dcpl_2831) , (and_dcpl_2832 & and_dcpl_2837) , (and_dcpl_2835
      & and_dcpl_2837) , (and_dcpl_2832 & and_dcpl_2843) , (and_dcpl_2835 & and_dcpl_2843)
      , (and_dcpl_2832 & and_dcpl_2849) , (and_dcpl_2835 & and_dcpl_2849) , ((else_7_if_1_div_9cyc_st_9[3])
      & (~ (else_7_if_1_div_9cyc_st_9[0])) & and_dcpl_2831) , and_2924_cse});
  assign mux1h_5_nl = MUX1HOT_v_13_10_2({(div_mgc_div_10_z[29:17]) , (div_mgc_div_11_z[29:17])
      , (div_mgc_div_12_z[29:17]) , (div_mgc_div_13_z[29:17]) , (div_mgc_div_14_z[29:17])
      , (div_mgc_div_15_z[29:17]) , (div_mgc_div_16_z[29:17]) , (div_mgc_div_17_z[29:17])
      , (div_mgc_div_18_z[29:17]) , (div_sdt_2_sva_duc[29:17])}, {and_2973_cse ,
      and_2976_cse , and_2979_cse , and_2982_cse , and_2985_cse , and_2988_cse ,
      and_2991_cse , and_2994_cse , and_2997_cse , and_3062_cse});
  assign nl_h_2_sva_1_sg1 = (mux1h_5_nl) + 13'b1;
  assign h_2_sva_1_sg1 = nl_h_2_sva_1_sg1[12:0];
  assign div_sdt_3_sva_duc_mx0 = MUX1HOT_v_30_10_2({(div_mgc_div_1_z[29:0]) , (div_mgc_div_2_z[29:0])
      , (div_mgc_div_3_z[29:0]) , (div_mgc_div_4_z[29:0]) , (div_mgc_div_5_z[29:0])
      , (div_mgc_div_6_z[29:0]) , (div_mgc_div_7_z[29:0]) , (div_mgc_div_8_z[29:0])
      , (div_mgc_div_9_z[29:0]) , div_sdt_3_sva_duc}, {and_3065_cse , and_3068_cse
      , and_3071_cse , and_3074_cse , and_3077_cse , and_3080_cse , and_3083_cse
      , and_3086_cse , and_3089_cse , and_3154_cse});
  assign h_2_lpi_dfm_1_sg2_1 = MUX1HOT_v_12_3_2({((div_sdt_3_sva_duc_mx0[29:18])
      + 12'b1) , (h_2_sva_1_sg1[12:1]) , (h_2_sva_duc_mx0[29:18])}, {else_7_nor_ssc
      , else_7_and_5_itm_9 , else_7_equal_svs_9});
  assign h_2_lpi_dfm_1_sg1_1 = MUX1HOT_s_1_3_2({(div_sdt_3_sva_duc_mx0[17]) , (h_2_sva_1_sg1[0])
      , (h_2_sva_duc_mx0[17])}, {else_7_nor_ssc , else_7_and_5_itm_9 , else_7_equal_svs_9});
  assign h_2_lpi_dfm_4 = MUX1HOT_v_17_12_2({(div_sdt_3_sva_duc_mx0[16:0]) , (div_mgc_div_10_z[16:0])
      , (div_mgc_div_11_z[16:0]) , (div_mgc_div_12_z[16:0]) , (div_mgc_div_13_z[16:0])
      , (div_mgc_div_14_z[16:0]) , (div_mgc_div_15_z[16:0]) , (div_mgc_div_16_z[16:0])
      , (div_mgc_div_17_z[16:0]) , (div_mgc_div_18_z[16:0]) , (div_sdt_2_sva_duc[16:0])
      , (h_2_sva_duc_mx0[16:0])}, {else_7_nor_ssc , (and_dcpl_2917 & and_dcpl_2915
      & else_7_and_5_itm_9) , (and_dcpl_2917 & and_dcpl_2914 & (else_7_else_1_if_div_9cyc_st_9[0])
      & else_7_and_5_itm_9) , (and_dcpl_2917 & and_dcpl_2924 & (~ (else_7_else_1_if_div_9cyc_st_9[0]))
      & else_7_and_5_itm_9) , (and_dcpl_2917 & and_dcpl_2924 & (else_7_else_1_if_div_9cyc_st_9[0])
      & else_7_and_5_itm_9) , (and_dcpl_2917 & and_dcpl_2934 & (~ (else_7_else_1_if_div_9cyc_st_9[0]))
      & else_7_and_5_itm_9) , (and_dcpl_2917 & and_dcpl_2934 & (else_7_else_1_if_div_9cyc_st_9[0])
      & else_7_and_5_itm_9) , (and_dcpl_2917 & and_dcpl_2944 & (~ (else_7_else_1_if_div_9cyc_st_9[0]))
      & else_7_and_5_itm_9) , (and_dcpl_2917 & and_dcpl_2944 & (else_7_else_1_if_div_9cyc_st_9[0])
      & else_7_and_5_itm_9) , (and_dcpl_2916 & (else_7_else_1_if_div_9cyc_st_9[3])
      & and_dcpl_2915 & else_7_and_5_itm_9) , ((and_3062_cse | or_dcpl_564) & else_7_and_5_itm_9)
      , else_7_equal_svs_9});
  assign else_7_nor_ssc = ~(else_7_else_1_equal_svs_st_9 | else_7_equal_svs_9);
  assign or_5023_cse = or_dcpl_857 | or_dcpl_855;
  assign or_5033_cse = or_dcpl_857 | or_dcpl_865;
  assign or_5043_cse = or_dcpl_877 | or_dcpl_855;
  assign or_5053_cse = or_dcpl_877 | or_dcpl_865;
  assign or_5063_cse = or_dcpl_857 | or_dcpl_895;
  assign or_5073_cse = or_dcpl_857 | or_dcpl_905;
  assign or_5083_cse = or_dcpl_877 | or_dcpl_895;
  assign or_5093_cse = or_dcpl_877 | or_dcpl_905;
  assign or_5103_cse = or_dcpl_857 | or_dcpl_935;
  assign or_5114_cse = or_dcpl_948 | or_dcpl_945;
  assign or_5126_cse = or_dcpl_948 | or_dcpl_957;
  assign or_5138_cse = or_dcpl_972 | or_dcpl_945;
  assign or_5150_cse = or_dcpl_972 | or_dcpl_957;
  assign or_5162_cse = or_dcpl_948 | or_dcpl_993;
  assign or_5174_cse = or_dcpl_948 | or_dcpl_1005;
  assign or_5186_cse = or_dcpl_972 | or_dcpl_993;
  assign or_5198_cse = or_dcpl_972 | or_dcpl_1005;
  assign or_5210_cse = or_dcpl_948 | or_dcpl_1041;
  assign or_5222_cse = or_dcpl_1056 | or_dcpl_1053;
  assign or_5234_cse = or_dcpl_1056 | or_dcpl_1065;
  assign or_5246_cse = or_dcpl_1080 | or_dcpl_1053;
  assign or_5258_cse = or_dcpl_1080 | or_dcpl_1065;
  assign else_7_equal_tmp = (r_sg1_lpi_dfm) == (mux1h_81_tmp);
  assign mux1h_81_tmp = MUX1HOT_v_16_3_2({(R_IN_rsc_mgc_in_wire_d[15:0]) , (B_IN_rsc_mgc_in_wire_d[15:0])
      , (G_IN_rsc_mgc_in_wire_d[15:0])}, {(~((if_if_acc_1_itm[17]) | (if_acc_itm[17])))
      , (((if_if_acc_1_itm[17]) & (~ (if_acc_itm[17]))) | ((else_1_if_acc_1_itm[17])
      & (if_acc_itm[17]))) , ((~ (else_1_if_acc_1_itm[17])) & (if_acc_itm[17]))});
  assign if_7_equal_tmp = (mux1h_81_tmp) == (min_sg1_lpi_dfm_3);
  assign nl_if_if_acc_1_itm = conv_s2u_17_18({(R_IN_rsc_mgc_in_wire_d[15:0]) , 1'b1})
      + conv_s2u_17_18({(~ (B_IN_rsc_mgc_in_wire_d[15:0])) , 1'b1});
  assign if_if_acc_1_itm = nl_if_if_acc_1_itm[17:0];
  assign nl_else_1_if_acc_1_itm = conv_s2u_17_18({(G_IN_rsc_mgc_in_wire_d[15:0])
      , 1'b1}) + conv_s2u_17_18({(~ (B_IN_rsc_mgc_in_wire_d[15:0])) , 1'b1});
  assign else_1_if_acc_1_itm = nl_else_1_if_acc_1_itm[17:0];
  assign nl_if_3_if_acc_1_itm = conv_s2u_17_18({(B_IN_rsc_mgc_in_wire_d[15:0]) ,
      1'b1}) + conv_s2u_17_18({(~ (R_IN_rsc_mgc_in_wire_d[15:0])) , 1'b1});
  assign if_3_if_acc_1_itm = nl_if_3_if_acc_1_itm[17:0];
  assign nl_else_5_if_acc_1_itm = conv_s2u_17_18({(B_IN_rsc_mgc_in_wire_d[15:0])
      , 1'b1}) + conv_s2u_17_18({(~ (G_IN_rsc_mgc_in_wire_d[15:0])) , 1'b1});
  assign else_5_if_acc_1_itm = nl_else_5_if_acc_1_itm[17:0];
  assign nl_else_7_acc_3_itm = ({mux1h_81_tmp , 1'b1}) + ({(~ min_sg1_lpi_dfm_3)
      , 1'b1});
  assign else_7_acc_3_itm = nl_else_7_acc_3_itm[16:0];
  assign nl_else_7_if_acc_tmp = conv_u2u_1_4(acc_5_itm[4]) + conv_u2u_3_4(acc_5_itm[3:1]);
  assign else_7_if_acc_tmp = nl_else_7_if_acc_tmp[3:0];
  assign nl_acc_5_itm = ({2'b10 , (else_7_if_acc_idiv[1:0]) , 1'b1}) + conv_u2s_4_5({(~
      (else_7_if_acc_idiv[2])) , 1'b1 , (~ (else_7_if_acc_idiv[2])) , (~ (else_7_if_acc_idiv[3]))});
  assign acc_5_itm = nl_acc_5_itm[4:0];
  assign nl_else_7_if_acc_idiv = else_7_if_div_9cyc + 4'b1;
  assign else_7_if_acc_idiv = nl_else_7_if_acc_idiv[3:0];
  assign nl_else_7_if_1_acc_1_itm = conv_s2u_17_18({g_sg1_lpi_dfm , 1'b1}) + conv_s2u_17_18({(~
      b_sg1_lpi_dfm) , 1'b1});
  assign else_7_if_1_acc_1_itm = nl_else_7_if_1_acc_1_itm[17:0];
  assign nl_else_7_if_1_acc_tmp = conv_u2u_1_4(acc_itm[4]) + conv_u2u_3_4(acc_itm[3:1]);
  assign else_7_if_1_acc_tmp = nl_else_7_if_1_acc_tmp[3:0];
  assign nl_acc_itm = ({2'b10 , (else_7_if_1_acc_idiv[1:0]) , 1'b1}) + conv_u2s_4_5({(~
      (else_7_if_1_acc_idiv[2])) , 1'b1 , (~ (else_7_if_1_acc_idiv[2])) , (~ (else_7_if_1_acc_idiv[3]))});
  assign acc_itm = nl_acc_itm[4:0];
  assign nl_else_7_if_1_acc_idiv = else_7_if_1_div_9cyc + 4'b1;
  assign else_7_if_1_acc_idiv = nl_else_7_if_1_acc_idiv[3:0];
  assign g_sg1_lpi_dfm = (G_IN_rsc_mgc_in_wire_d[15:0]) & ({{15{unequal_tmp}}, unequal_tmp});
  assign b_sg1_lpi_dfm = (B_IN_rsc_mgc_in_wire_d[15:0]) & ({{15{unequal_tmp}}, unequal_tmp});
  assign nl_else_7_else_1_if_acc_2_itm = conv_s2u_17_18({b_sg1_lpi_dfm , 1'b1}) +
      conv_s2u_17_18({(~ r_sg1_lpi_dfm) , 1'b1});
  assign else_7_else_1_if_acc_2_itm = nl_else_7_else_1_if_acc_2_itm[17:0];
  assign nl_else_7_else_1_if_acc_tmp = conv_u2u_1_4(acc_6_itm[4]) + conv_u2u_3_4(acc_6_itm[3:1]);
  assign else_7_else_1_if_acc_tmp = nl_else_7_else_1_if_acc_tmp[3:0];
  assign nl_acc_6_itm = ({2'b10 , (else_7_else_1_if_acc_idiv[1:0]) , 1'b1}) + conv_u2s_4_5({(~
      (else_7_else_1_if_acc_idiv[2])) , 1'b1 , (~ (else_7_else_1_if_acc_idiv[2]))
      , (~ (else_7_else_1_if_acc_idiv[3]))});
  assign acc_6_itm = nl_acc_6_itm[4:0];
  assign nl_else_7_else_1_if_acc_idiv = else_7_else_1_if_div_9cyc + 4'b1;
  assign else_7_else_1_if_acc_idiv = nl_else_7_else_1_if_acc_idiv[3:0];
  assign r_sg1_lpi_dfm = (R_IN_rsc_mgc_in_wire_d[15:0]) & ({{15{unequal_tmp}}, unequal_tmp});
  assign nl_else_7_else_1_else_acc_2_itm = conv_s2u_17_18({r_sg1_lpi_dfm , 1'b1})
      + conv_s2u_17_18({(~ g_sg1_lpi_dfm) , 1'b1});
  assign else_7_else_1_else_acc_2_itm = nl_else_7_else_1_else_acc_2_itm[17:0];
  assign nl_else_7_else_1_else_acc_tmp = conv_u2u_1_4(acc_7_itm[4]) + conv_u2u_3_4(acc_7_itm[3:1]);
  assign else_7_else_1_else_acc_tmp = nl_else_7_else_1_else_acc_tmp[3:0];
  assign nl_acc_7_itm = ({2'b10 , (else_7_else_1_else_acc_idiv[1:0]) , 1'b1}) + conv_u2s_4_5({(~
      (else_7_else_1_else_acc_idiv[2])) , 1'b1 , (~ (else_7_else_1_else_acc_idiv[2]))
      , (~ (else_7_else_1_else_acc_idiv[3]))});
  assign acc_7_itm = nl_acc_7_itm[4:0];
  assign nl_else_7_else_1_else_acc_idiv = else_7_else_1_else_div_9cyc + 4'b1;
  assign else_7_else_1_else_acc_idiv = nl_else_7_else_1_else_acc_idiv[3:0];
  assign else_7_else_1_equal_tmp = (g_sg1_lpi_dfm) == (mux1h_81_tmp);
  assign unequal_tmp = (mux1h_81_tmp[15]) | (mux1h_81_tmp[14]) | (mux1h_81_tmp[13])
      | (mux1h_81_tmp[12]) | (mux1h_81_tmp[11]) | (mux1h_81_tmp[10]) | (mux1h_81_tmp[9])
      | (mux1h_81_tmp[8]) | (mux1h_81_tmp[7]) | (mux1h_81_tmp[6]) | (mux1h_81_tmp[5])
      | (mux1h_81_tmp[4]) | (mux1h_81_tmp[3]) | (mux1h_81_tmp[2]) | (mux1h_81_tmp[1])
      | (mux1h_81_tmp[0]);
  assign min_sg1_lpi_dfm_3 = MUX1HOT_v_16_3_2({(R_IN_rsc_mgc_in_wire_d[15:0]) , (B_IN_rsc_mgc_in_wire_d[15:0])
      , (G_IN_rsc_mgc_in_wire_d[15:0])}, {(~((if_3_if_acc_1_itm[17]) | (if_3_acc_itm[17])))
      , (((if_3_if_acc_1_itm[17]) & (~ (if_3_acc_itm[17]))) | ((else_5_if_acc_1_itm[17])
      & (if_3_acc_itm[17]))) , ((~ (else_5_if_acc_1_itm[17])) & (if_3_acc_itm[17]))});
  assign nl_if_3_acc_itm = conv_s2u_17_18({(G_IN_rsc_mgc_in_wire_d[15:0]) , 1'b1})
      + conv_s2u_17_18({(~ (R_IN_rsc_mgc_in_wire_d[15:0])) , 1'b1});
  assign if_3_acc_itm = nl_if_3_acc_itm[17:0];
  assign nl_if_acc_itm = conv_s2u_17_18({(R_IN_rsc_mgc_in_wire_d[15:0]) , 1'b1})
      + conv_s2u_17_18({(~ (G_IN_rsc_mgc_in_wire_d[15:0])) , 1'b1});
  assign if_acc_itm = nl_if_acc_itm[17:0];
  assign and_dcpl_15 = ~((else_7_if_div_9cyc_st_7[3]) | (else_7_if_div_9cyc_st_7[0]));
  assign and_dcpl_17 = (~ if_7_equal_svs_st_7) & main_stage_0_8;
  assign and_dcpl_27 = (~ (else_7_if_div_9cyc_st_7[3])) & (else_7_if_div_9cyc_st_7[0]);
  assign and_dcpl_124 = ~((else_7_if_1_div_9cyc_st_7[3]) | (else_7_if_1_div_9cyc_st_7[0]));
  assign and_dcpl_136 = (~ (else_7_if_1_div_9cyc_st_7[3])) & (else_7_if_1_div_9cyc_st_7[0]);
  assign and_dcpl_234 = ~((else_7_else_1_if_div_9cyc_st_7[0]) | (else_7_else_1_if_div_9cyc_st_7[1]));
  assign and_dcpl_235 = ~((else_7_else_1_if_div_9cyc_st_7[2]) | (else_7_else_1_if_div_9cyc_st_7[3]));
  assign and_dcpl_248 = (else_7_else_1_if_div_9cyc_st_7[0]) & (~ (else_7_else_1_if_div_9cyc_st_7[1]));
  assign and_dcpl_262 = (~ (else_7_else_1_if_div_9cyc_st_7[0])) & (else_7_else_1_if_div_9cyc_st_7[1]);
  assign and_dcpl_276 = (else_7_else_1_if_div_9cyc_st_7[0]) & (else_7_else_1_if_div_9cyc_st_7[1]);
  assign and_dcpl_291 = (else_7_else_1_if_div_9cyc_st_7[2]) & (~ (else_7_else_1_if_div_9cyc_st_7[3]));
  assign and_dcpl_363 = ~((else_7_else_1_else_div_9cyc_st_7[0]) | (else_7_else_1_else_div_9cyc_st_7[1]));
  assign and_dcpl_364 = ~((else_7_else_1_else_div_9cyc_st_7[2]) | (else_7_else_1_else_div_9cyc_st_7[3]));
  assign and_dcpl_377 = (else_7_else_1_else_div_9cyc_st_7[0]) & (~ (else_7_else_1_else_div_9cyc_st_7[1]));
  assign and_dcpl_391 = (~ (else_7_else_1_else_div_9cyc_st_7[0])) & (else_7_else_1_else_div_9cyc_st_7[1]);
  assign and_dcpl_405 = (else_7_else_1_else_div_9cyc_st_7[0]) & (else_7_else_1_else_div_9cyc_st_7[1]);
  assign and_dcpl_420 = (else_7_else_1_else_div_9cyc_st_7[2]) & (~ (else_7_else_1_else_div_9cyc_st_7[3]));
  assign and_506_cse = (~ if_7_equal_svs_st_6) & main_stage_0_7;
  assign and_dcpl_496 = ~((else_7_if_1_div_9cyc_st_6[3]) | (else_7_if_1_div_9cyc_st_6[0]));
  assign and_dcpl_508 = (~ (else_7_if_1_div_9cyc_st_6[3])) & (else_7_if_1_div_9cyc_st_6[0]);
  assign and_dcpl_606 = ~((else_7_else_1_if_div_9cyc_st_6[0]) | (else_7_else_1_if_div_9cyc_st_6[1]));
  assign and_dcpl_607 = ~((else_7_else_1_if_div_9cyc_st_6[2]) | (else_7_else_1_if_div_9cyc_st_6[3]));
  assign and_dcpl_620 = (else_7_else_1_if_div_9cyc_st_6[0]) & (~ (else_7_else_1_if_div_9cyc_st_6[1]));
  assign and_dcpl_634 = (~ (else_7_else_1_if_div_9cyc_st_6[0])) & (else_7_else_1_if_div_9cyc_st_6[1]);
  assign and_dcpl_648 = (else_7_else_1_if_div_9cyc_st_6[0]) & (else_7_else_1_if_div_9cyc_st_6[1]);
  assign and_dcpl_663 = (else_7_else_1_if_div_9cyc_st_6[2]) & (~ (else_7_else_1_if_div_9cyc_st_6[3]));
  assign and_dcpl_735 = ~((else_7_else_1_else_div_9cyc_st_6[0]) | (else_7_else_1_else_div_9cyc_st_6[1]));
  assign and_dcpl_736 = ~((else_7_else_1_else_div_9cyc_st_6[2]) | (else_7_else_1_else_div_9cyc_st_6[3]));
  assign and_dcpl_749 = (else_7_else_1_else_div_9cyc_st_6[0]) & (~ (else_7_else_1_else_div_9cyc_st_6[1]));
  assign and_dcpl_763 = (~ (else_7_else_1_else_div_9cyc_st_6[0])) & (else_7_else_1_else_div_9cyc_st_6[1]);
  assign and_dcpl_777 = (else_7_else_1_else_div_9cyc_st_6[0]) & (else_7_else_1_else_div_9cyc_st_6[1]);
  assign and_dcpl_792 = (else_7_else_1_else_div_9cyc_st_6[2]) & (~ (else_7_else_1_else_div_9cyc_st_6[3]));
  assign and_878_cse = (~ if_7_equal_svs_st_5) & main_stage_0_6;
  assign and_dcpl_868 = ~((else_7_if_1_div_9cyc_st_5[1]) | (else_7_if_1_div_9cyc_st_5[2]));
  assign and_dcpl_892 = (else_7_if_1_div_9cyc_st_5[1]) & (~ (else_7_if_1_div_9cyc_st_5[2]));
  assign and_dcpl_916 = (~ (else_7_if_1_div_9cyc_st_5[1])) & (else_7_if_1_div_9cyc_st_5[2]);
  assign and_dcpl_940 = (else_7_if_1_div_9cyc_st_5[1]) & (else_7_if_1_div_9cyc_st_5[2]);
  assign and_dcpl_978 = ~((else_7_else_1_if_div_9cyc_st_5[0]) | (else_7_else_1_if_div_9cyc_st_5[1]));
  assign and_dcpl_979 = ~((else_7_else_1_if_div_9cyc_st_5[2]) | (else_7_else_1_if_div_9cyc_st_5[3]));
  assign and_dcpl_992 = (else_7_else_1_if_div_9cyc_st_5[0]) & (~ (else_7_else_1_if_div_9cyc_st_5[1]));
  assign and_dcpl_1006 = (~ (else_7_else_1_if_div_9cyc_st_5[0])) & (else_7_else_1_if_div_9cyc_st_5[1]);
  assign and_dcpl_1020 = (else_7_else_1_if_div_9cyc_st_5[0]) & (else_7_else_1_if_div_9cyc_st_5[1]);
  assign and_dcpl_1035 = (else_7_else_1_if_div_9cyc_st_5[2]) & (~ (else_7_else_1_if_div_9cyc_st_5[3]));
  assign and_dcpl_1107 = ~((else_7_else_1_else_div_9cyc_st_5[0]) | (else_7_else_1_else_div_9cyc_st_5[1]));
  assign and_dcpl_1108 = ~((else_7_else_1_else_div_9cyc_st_5[2]) | (else_7_else_1_else_div_9cyc_st_5[3]));
  assign and_dcpl_1121 = (else_7_else_1_else_div_9cyc_st_5[0]) & (~ (else_7_else_1_else_div_9cyc_st_5[1]));
  assign and_dcpl_1135 = (~ (else_7_else_1_else_div_9cyc_st_5[0])) & (else_7_else_1_else_div_9cyc_st_5[1]);
  assign and_dcpl_1149 = (else_7_else_1_else_div_9cyc_st_5[0]) & (else_7_else_1_else_div_9cyc_st_5[1]);
  assign and_dcpl_1164 = (else_7_else_1_else_div_9cyc_st_5[2]) & (~ (else_7_else_1_else_div_9cyc_st_5[3]));
  assign and_1250_cse = (~ if_7_equal_svs_st_4) & main_stage_0_5;
  assign and_dcpl_1240 = ~((else_7_if_1_div_9cyc_st_4[3]) | (else_7_if_1_div_9cyc_st_4[0]));
  assign and_dcpl_1252 = (~ (else_7_if_1_div_9cyc_st_4[3])) & (else_7_if_1_div_9cyc_st_4[0]);
  assign and_dcpl_1350 = ~((else_7_else_1_if_div_9cyc_st_4[0]) | (else_7_else_1_if_div_9cyc_st_4[1]));
  assign and_dcpl_1351 = ~((else_7_else_1_if_div_9cyc_st_4[2]) | (else_7_else_1_if_div_9cyc_st_4[3]));
  assign and_dcpl_1364 = (else_7_else_1_if_div_9cyc_st_4[0]) & (~ (else_7_else_1_if_div_9cyc_st_4[1]));
  assign and_dcpl_1378 = (~ (else_7_else_1_if_div_9cyc_st_4[0])) & (else_7_else_1_if_div_9cyc_st_4[1]);
  assign and_dcpl_1392 = (else_7_else_1_if_div_9cyc_st_4[0]) & (else_7_else_1_if_div_9cyc_st_4[1]);
  assign and_dcpl_1407 = (else_7_else_1_if_div_9cyc_st_4[2]) & (~ (else_7_else_1_if_div_9cyc_st_4[3]));
  assign and_dcpl_1479 = ~((else_7_else_1_else_div_9cyc_st_4[0]) | (else_7_else_1_else_div_9cyc_st_4[1]));
  assign and_dcpl_1480 = ~((else_7_else_1_else_div_9cyc_st_4[2]) | (else_7_else_1_else_div_9cyc_st_4[3]));
  assign and_dcpl_1493 = (else_7_else_1_else_div_9cyc_st_4[0]) & (~ (else_7_else_1_else_div_9cyc_st_4[1]));
  assign and_dcpl_1507 = (~ (else_7_else_1_else_div_9cyc_st_4[0])) & (else_7_else_1_else_div_9cyc_st_4[1]);
  assign and_dcpl_1521 = (else_7_else_1_else_div_9cyc_st_4[0]) & (else_7_else_1_else_div_9cyc_st_4[1]);
  assign and_dcpl_1536 = (else_7_else_1_else_div_9cyc_st_4[2]) & (~ (else_7_else_1_else_div_9cyc_st_4[3]));
  assign and_1622_cse = (~ if_7_equal_svs_st_3) & main_stage_0_4;
  assign and_dcpl_1612 = ~((else_7_if_1_div_9cyc_st_3[3]) | (else_7_if_1_div_9cyc_st_3[1]));
  assign and_dcpl_1636 = (~ (else_7_if_1_div_9cyc_st_3[3])) & (else_7_if_1_div_9cyc_st_3[1]);
  assign and_dcpl_1722 = ~((else_7_else_1_if_div_9cyc_st_3[1]) | (else_7_else_1_if_div_9cyc_st_3[2]));
  assign and_dcpl_1723 = ~((else_7_else_1_if_div_9cyc_st_3[0]) | (else_7_else_1_if_div_9cyc_st_3[3]));
  assign and_dcpl_1737 = (else_7_else_1_if_div_9cyc_st_3[0]) & (~ (else_7_else_1_if_div_9cyc_st_3[3]));
  assign and_dcpl_1750 = (else_7_else_1_if_div_9cyc_st_3[1]) & (~ (else_7_else_1_if_div_9cyc_st_3[2]));
  assign and_dcpl_1778 = (~ (else_7_else_1_if_div_9cyc_st_3[1])) & (else_7_else_1_if_div_9cyc_st_3[2]);
  assign and_dcpl_1806 = (else_7_else_1_if_div_9cyc_st_3[1]) & (else_7_else_1_if_div_9cyc_st_3[2]);
  assign and_dcpl_1851 = ~((else_7_else_1_else_div_9cyc_st_3[0]) | (else_7_else_1_else_div_9cyc_st_3[1]));
  assign and_dcpl_1852 = ~((else_7_else_1_else_div_9cyc_st_3[2]) | (else_7_else_1_else_div_9cyc_st_3[3]));
  assign and_dcpl_1865 = (else_7_else_1_else_div_9cyc_st_3[0]) & (~ (else_7_else_1_else_div_9cyc_st_3[1]));
  assign and_dcpl_1879 = (~ (else_7_else_1_else_div_9cyc_st_3[0])) & (else_7_else_1_else_div_9cyc_st_3[1]);
  assign and_dcpl_1893 = (else_7_else_1_else_div_9cyc_st_3[0]) & (else_7_else_1_else_div_9cyc_st_3[1]);
  assign and_dcpl_1908 = (else_7_else_1_else_div_9cyc_st_3[2]) & (~ (else_7_else_1_else_div_9cyc_st_3[3]));
  assign and_1994_cse = main_stage_0_3 & (~ if_7_equal_svs_st_2);
  assign and_dcpl_1984 = ~((else_7_if_1_div_9cyc_st_2[3]) | (else_7_if_1_div_9cyc_st_2[1]));
  assign and_dcpl_2008 = (~ (else_7_if_1_div_9cyc_st_2[3])) & (else_7_if_1_div_9cyc_st_2[1]);
  assign and_dcpl_2094 = ~((else_7_else_1_if_div_9cyc_st_2[2]) | (else_7_else_1_if_div_9cyc_st_2[0]));
  assign and_dcpl_2095 = ~((else_7_else_1_if_div_9cyc_st_2[3]) | (else_7_else_1_if_div_9cyc_st_2[1]));
  assign and_dcpl_2108 = (~ (else_7_else_1_if_div_9cyc_st_2[2])) & (else_7_else_1_if_div_9cyc_st_2[0]);
  assign and_dcpl_2123 = (~ (else_7_else_1_if_div_9cyc_st_2[3])) & (else_7_else_1_if_div_9cyc_st_2[1]);
  assign and_dcpl_2150 = (else_7_else_1_if_div_9cyc_st_2[2]) & (~ (else_7_else_1_if_div_9cyc_st_2[0]));
  assign and_dcpl_2164 = (else_7_else_1_if_div_9cyc_st_2[2]) & (else_7_else_1_if_div_9cyc_st_2[0]);
  assign and_dcpl_2223 = ~((else_7_else_1_else_div_9cyc_st_2[1]) | (else_7_else_1_else_div_9cyc_st_2[0]));
  assign and_dcpl_2224 = ~((else_7_else_1_else_div_9cyc_st_2[2]) | (else_7_else_1_else_div_9cyc_st_2[3]));
  assign and_dcpl_2237 = (~ (else_7_else_1_else_div_9cyc_st_2[1])) & (else_7_else_1_else_div_9cyc_st_2[0]);
  assign and_dcpl_2251 = (else_7_else_1_else_div_9cyc_st_2[1]) & (~ (else_7_else_1_else_div_9cyc_st_2[0]));
  assign and_dcpl_2265 = (else_7_else_1_else_div_9cyc_st_2[1]) & (else_7_else_1_else_div_9cyc_st_2[0]);
  assign and_dcpl_2280 = (else_7_else_1_else_div_9cyc_st_2[2]) & (~ (else_7_else_1_else_div_9cyc_st_2[3]));
  assign and_2366_cse = (~ if_7_equal_svs_st_1) & main_stage_0_2;
  assign and_dcpl_2356 = ~((else_7_if_1_div_9cyc[3]) | (else_7_if_1_div_9cyc[1]));
  assign and_dcpl_2380 = (~ (else_7_if_1_div_9cyc[3])) & (else_7_if_1_div_9cyc[1]);
  assign and_dcpl_2741 = ~((else_7_if_div_9cyc_st_9[1]) | (else_7_if_div_9cyc_st_9[2]));
  assign and_dcpl_2742 = ~((else_7_if_div_9cyc_st_9[3]) | (else_7_if_div_9cyc_st_9[0]));
  assign and_dcpl_2746 = (~ (else_7_if_div_9cyc_st_9[3])) & (else_7_if_div_9cyc_st_9[0]);
  assign and_dcpl_2749 = (else_7_if_div_9cyc_st_9[1]) & (~ (else_7_if_div_9cyc_st_9[2]));
  assign and_dcpl_2757 = (~ (else_7_if_div_9cyc_st_9[1])) & (else_7_if_div_9cyc_st_9[2]);
  assign and_dcpl_2765 = (else_7_if_div_9cyc_st_9[1]) & (else_7_if_div_9cyc_st_9[2]);
  assign or_tmp_4 = (((else_7_if_div_9cyc_st_9[2]) | (else_7_if_div_9cyc_st_9[1])
      | (else_7_if_div_9cyc_st_9[0])) & (else_7_if_div_9cyc_st_9[3])) | (~((max_sg1_lpi_dfm_3_st_9[0])
      | (max_sg1_lpi_dfm_3_st_9[1]) | (max_sg1_lpi_dfm_3_st_9[2]) | (max_sg1_lpi_dfm_3_st_9[3])
      | (max_sg1_lpi_dfm_3_st_9[4]) | (max_sg1_lpi_dfm_3_st_9[5]) | (max_sg1_lpi_dfm_3_st_9[6])
      | (max_sg1_lpi_dfm_3_st_9[7]) | (max_sg1_lpi_dfm_3_st_9[8]) | (max_sg1_lpi_dfm_3_st_9[9])
      | (max_sg1_lpi_dfm_3_st_9[10]) | (max_sg1_lpi_dfm_3_st_9[11]) | (max_sg1_lpi_dfm_3_st_9[12])
      | (max_sg1_lpi_dfm_3_st_9[13]) | (max_sg1_lpi_dfm_3_st_9[14]) | (max_sg1_lpi_dfm_3_st_9[15])));
  assign and_dcpl_2777 = ~((else_7_if_div_9cyc_st_9[0]) | (else_7_if_div_9cyc_st_9[1]));
  assign and_dcpl_2778 = and_dcpl_2777 & (~ (else_7_if_div_9cyc_st_9[2]));
  assign and_dcpl_2780 = and_9092_cse & (~ (else_7_if_div_9cyc_st_9[3]));
  assign and_dcpl_2783 = (else_7_if_div_9cyc_st_9[0]) & (~ (else_7_if_div_9cyc_st_9[1]));
  assign and_dcpl_2789 = (~ (else_7_if_div_9cyc_st_9[0])) & (else_7_if_div_9cyc_st_9[1]);
  assign and_dcpl_2795 = (else_7_if_div_9cyc_st_9[0]) & (else_7_if_div_9cyc_st_9[1]);
  assign or_dcpl_555 = if_7_equal_svs_9 | (~ main_stage_0_10);
  assign and_dcpl_2831 = ~((else_7_if_1_div_9cyc_st_9[1]) | (else_7_if_1_div_9cyc_st_9[2]));
  assign and_dcpl_2832 = ~((else_7_if_1_div_9cyc_st_9[3]) | (else_7_if_1_div_9cyc_st_9[0]));
  assign and_dcpl_2835 = (~ (else_7_if_1_div_9cyc_st_9[3])) & (else_7_if_1_div_9cyc_st_9[0]);
  assign and_dcpl_2837 = (else_7_if_1_div_9cyc_st_9[1]) & (~ (else_7_if_1_div_9cyc_st_9[2]));
  assign and_dcpl_2843 = (~ (else_7_if_1_div_9cyc_st_9[1])) & (else_7_if_1_div_9cyc_st_9[2]);
  assign and_dcpl_2849 = (else_7_if_1_div_9cyc_st_9[1]) & (else_7_if_1_div_9cyc_st_9[2]);
  assign and_dcpl_2859 = ~((else_7_if_1_div_9cyc_st_9[0]) | (else_7_if_1_div_9cyc_st_9[1]));
  assign and_dcpl_2860 = and_dcpl_2859 & (~ (else_7_if_1_div_9cyc_st_9[2]));
  assign and_dcpl_2863 = and_9092_cse & else_7_equal_svs_9 & (~ (else_7_if_1_div_9cyc_st_9[3]));
  assign and_dcpl_2865 = (else_7_if_1_div_9cyc_st_9[0]) & (~ (else_7_if_1_div_9cyc_st_9[1]));
  assign and_dcpl_2871 = (~ (else_7_if_1_div_9cyc_st_9[0])) & (else_7_if_1_div_9cyc_st_9[1]);
  assign and_dcpl_2877 = (else_7_if_1_div_9cyc_st_9[0]) & (else_7_if_1_div_9cyc_st_9[1]);
  assign and_dcpl_2914 = ~((else_7_else_1_if_div_9cyc_st_9[2]) | (else_7_else_1_if_div_9cyc_st_9[1]));
  assign and_dcpl_2915 = and_dcpl_2914 & (~ (else_7_else_1_if_div_9cyc_st_9[0]));
  assign and_dcpl_2916 = (~ else_7_equal_svs_9) & else_7_else_1_equal_svs_st_9;
  assign and_dcpl_2917 = and_dcpl_2916 & (~ (else_7_else_1_if_div_9cyc_st_9[3]));
  assign and_dcpl_2924 = (~ (else_7_else_1_if_div_9cyc_st_9[2])) & (else_7_else_1_if_div_9cyc_st_9[1]);
  assign and_dcpl_2934 = (else_7_else_1_if_div_9cyc_st_9[2]) & (~ (else_7_else_1_if_div_9cyc_st_9[1]));
  assign and_dcpl_2944 = (else_7_else_1_if_div_9cyc_st_9[2]) & (else_7_else_1_if_div_9cyc_st_9[1]);
  assign or_dcpl_564 = else_7_equal_svs_9 | (~ else_7_else_1_equal_svs_st_9);
  assign and_dcpl_2960 = ~((else_7_else_1_if_div_9cyc_st_9[1]) | (else_7_else_1_if_div_9cyc_st_9[0]));
  assign and_dcpl_2961 = ~((else_7_else_1_if_div_9cyc_st_9[3]) | (else_7_else_1_if_div_9cyc_st_9[2]));
  assign and_2973_cse = and_dcpl_2961 & and_dcpl_2960;
  assign and_dcpl_2963 = (~ (else_7_else_1_if_div_9cyc_st_9[1])) & (else_7_else_1_if_div_9cyc_st_9[0]);
  assign and_2976_cse = and_dcpl_2961 & and_dcpl_2963;
  assign and_dcpl_2966 = (else_7_else_1_if_div_9cyc_st_9[1]) & (~ (else_7_else_1_if_div_9cyc_st_9[0]));
  assign and_2979_cse = and_dcpl_2961 & and_dcpl_2966;
  assign and_dcpl_2969 = (else_7_else_1_if_div_9cyc_st_9[1]) & (else_7_else_1_if_div_9cyc_st_9[0]);
  assign and_2982_cse = and_dcpl_2961 & and_dcpl_2969;
  assign and_dcpl_2973 = (~ (else_7_else_1_if_div_9cyc_st_9[3])) & (else_7_else_1_if_div_9cyc_st_9[2]);
  assign and_2985_cse = and_dcpl_2973 & and_dcpl_2960;
  assign and_2988_cse = and_dcpl_2973 & and_dcpl_2963;
  assign and_2991_cse = and_dcpl_2973 & and_dcpl_2966;
  assign and_2994_cse = and_dcpl_2973 & and_dcpl_2969;
  assign and_2997_cse = (else_7_else_1_if_div_9cyc_st_9[3]) & (~ (else_7_else_1_if_div_9cyc_st_9[2]))
      & and_dcpl_2960;
  assign and_dcpl_2993 = and_9092_cse & and_dcpl_2916;
  assign and_dcpl_3052 = ~((else_7_else_1_else_div_9cyc_st_9[1]) | (else_7_else_1_else_div_9cyc_st_9[2]));
  assign and_dcpl_3053 = ~((else_7_else_1_else_div_9cyc_st_9[3]) | (else_7_else_1_else_div_9cyc_st_9[0]));
  assign and_3065_cse = and_dcpl_3053 & and_dcpl_3052;
  assign and_dcpl_3056 = (~ (else_7_else_1_else_div_9cyc_st_9[3])) & (else_7_else_1_else_div_9cyc_st_9[0]);
  assign and_3068_cse = and_dcpl_3056 & and_dcpl_3052;
  assign and_dcpl_3058 = (else_7_else_1_else_div_9cyc_st_9[1]) & (~ (else_7_else_1_else_div_9cyc_st_9[2]));
  assign and_3071_cse = and_dcpl_3053 & and_dcpl_3058;
  assign and_3074_cse = and_dcpl_3056 & and_dcpl_3058;
  assign and_dcpl_3064 = (~ (else_7_else_1_else_div_9cyc_st_9[1])) & (else_7_else_1_else_div_9cyc_st_9[2]);
  assign and_3077_cse = and_dcpl_3053 & and_dcpl_3064;
  assign and_3080_cse = and_dcpl_3056 & and_dcpl_3064;
  assign and_dcpl_3070 = (else_7_else_1_else_div_9cyc_st_9[1]) & (else_7_else_1_else_div_9cyc_st_9[2]);
  assign and_3083_cse = and_dcpl_3053 & and_dcpl_3070;
  assign and_3086_cse = and_dcpl_3056 & and_dcpl_3070;
  assign and_3089_cse = (else_7_else_1_else_div_9cyc_st_9[3]) & (~ (else_7_else_1_else_div_9cyc_st_9[0]))
      & and_dcpl_3052;
  assign and_dcpl_3085 = and_9092_cse & (~(else_7_equal_svs_9 | else_7_else_1_equal_svs_st_9));
  assign and_dcpl_3144 = ~((else_7_if_acc_tmp[1]) | (else_7_if_acc_tmp[0]));
  assign and_dcpl_3145 = ~(if_7_equal_tmp | (else_7_if_acc_tmp[3]));
  assign and_dcpl_3146 = and_dcpl_3145 & (~ (else_7_if_acc_tmp[2]));
  assign and_dcpl_3149 = ~((else_7_if_div_9cyc_st_1[2]) | (else_7_if_div_9cyc_st_1[1]));
  assign and_dcpl_3150 = and_dcpl_3149 & (~ (else_7_if_div_9cyc_st_1[0]));
  assign and_dcpl_3152 = and_2366_cse & (~ (else_7_if_div_9cyc_st_1[3]));
  assign or_tmp_6 = (max_sg1_lpi_dfm_3_st_1[0]) | (max_sg1_lpi_dfm_3_st_1[15]) |
      (max_sg1_lpi_dfm_3_st_1[14]) | (max_sg1_lpi_dfm_3_st_1[13]) | (max_sg1_lpi_dfm_3_st_1[12])
      | (max_sg1_lpi_dfm_3_st_1[11]) | (max_sg1_lpi_dfm_3_st_1[10]) | (max_sg1_lpi_dfm_3_st_1[9])
      | (max_sg1_lpi_dfm_3_st_1[8]) | (max_sg1_lpi_dfm_3_st_1[7]) | (max_sg1_lpi_dfm_3_st_1[6])
      | (max_sg1_lpi_dfm_3_st_1[5]) | (max_sg1_lpi_dfm_3_st_1[4]) | (max_sg1_lpi_dfm_3_st_1[3])
      | (max_sg1_lpi_dfm_3_st_1[2]) | (max_sg1_lpi_dfm_3_st_1[1]);
  assign or_tmp_7 = (mux1h_81_tmp[15]) | (mux1h_81_tmp[14]) | (mux1h_81_tmp[13])
      | (mux1h_81_tmp[12]) | (mux1h_81_tmp[11]) | (mux1h_81_tmp[10]) | (mux1h_81_tmp[9])
      | (mux1h_81_tmp[8]) | (mux1h_81_tmp[7]) | (mux1h_81_tmp[6]) | (mux1h_81_tmp[5])
      | (mux1h_81_tmp[4]) | (mux1h_81_tmp[3]) | (mux1h_81_tmp[2]) | (mux1h_81_tmp[1])
      | (mux1h_81_tmp[0]);
  assign not_tmp_146 = ~(or_tmp_7 | (~ or_tmp_6));
  assign and_dcpl_3155 = ~((else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[1]));
  assign and_dcpl_3156 = and_dcpl_3155 & (~ (else_7_if_div_9cyc_st_2[2]));
  assign and_dcpl_3158 = and_1994_cse & (~ (else_7_if_div_9cyc_st_2[3]));
  assign or_tmp_9 = (else_7_if_acc_tmp[3]) | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[1])
      | (else_7_if_acc_tmp[0]) | if_7_equal_tmp;
  assign or_tmp_10 = (max_sg1_lpi_dfm_3_st_1[0]) | (max_sg1_lpi_dfm_3_st_1[1]) |
      (max_sg1_lpi_dfm_3_st_1[2]) | (max_sg1_lpi_dfm_3_st_1[3]) | (max_sg1_lpi_dfm_3_st_1[4])
      | (max_sg1_lpi_dfm_3_st_1[5]) | (max_sg1_lpi_dfm_3_st_1[6]) | (max_sg1_lpi_dfm_3_st_1[7])
      | (max_sg1_lpi_dfm_3_st_1[8]) | (max_sg1_lpi_dfm_3_st_1[9]) | (max_sg1_lpi_dfm_3_st_1[10])
      | (max_sg1_lpi_dfm_3_st_1[11]) | (max_sg1_lpi_dfm_3_st_1[12]) | (max_sg1_lpi_dfm_3_st_1[13])
      | (max_sg1_lpi_dfm_3_st_1[14]) | (max_sg1_lpi_dfm_3_st_1[15]);
  assign or_tmp_12 = (max_sg1_lpi_dfm_3_st_2[0]) | (max_sg1_lpi_dfm_3_st_2[1]) |
      (max_sg1_lpi_dfm_3_st_2[2]) | (max_sg1_lpi_dfm_3_st_2[3]) | (max_sg1_lpi_dfm_3_st_2[4])
      | (max_sg1_lpi_dfm_3_st_2[5]) | (max_sg1_lpi_dfm_3_st_2[6]) | (max_sg1_lpi_dfm_3_st_2[7])
      | (max_sg1_lpi_dfm_3_st_2[8]) | (max_sg1_lpi_dfm_3_st_2[9]) | (max_sg1_lpi_dfm_3_st_2[10])
      | (max_sg1_lpi_dfm_3_st_2[11]) | (max_sg1_lpi_dfm_3_st_2[12]) | (max_sg1_lpi_dfm_3_st_2[13])
      | (max_sg1_lpi_dfm_3_st_2[14]) | (max_sg1_lpi_dfm_3_st_2[15]);
  assign or_612_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (else_7_if_div_9cyc_st_1[0]) | (else_7_if_div_9cyc_st_1[1]) | (else_7_if_div_9cyc_st_1[2])
      | (else_7_if_div_9cyc_st_1[3]);
  assign and_tmp = or_612_cse & or_tmp_12;
  assign and_dcpl_3161 = ~((else_7_if_div_9cyc_st_3[1]) | (else_7_if_div_9cyc_st_3[2]));
  assign and_dcpl_3162 = and_dcpl_3161 & (~ (else_7_if_div_9cyc_st_3[3]));
  assign and_dcpl_3164 = and_1622_cse & (~ (else_7_if_div_9cyc_st_3[0]));
  assign or_tmp_15 = (max_sg1_lpi_dfm_3_st_3[0]) | (max_sg1_lpi_dfm_3_st_3[1]) |
      (max_sg1_lpi_dfm_3_st_3[2]) | (max_sg1_lpi_dfm_3_st_3[3]) | (max_sg1_lpi_dfm_3_st_3[4])
      | (max_sg1_lpi_dfm_3_st_3[5]) | (max_sg1_lpi_dfm_3_st_3[6]) | (max_sg1_lpi_dfm_3_st_3[7])
      | (max_sg1_lpi_dfm_3_st_3[8]) | (max_sg1_lpi_dfm_3_st_3[9]) | (max_sg1_lpi_dfm_3_st_3[10])
      | (max_sg1_lpi_dfm_3_st_3[11]) | (max_sg1_lpi_dfm_3_st_3[12]) | (max_sg1_lpi_dfm_3_st_3[13])
      | (max_sg1_lpi_dfm_3_st_3[14]) | (max_sg1_lpi_dfm_3_st_3[15]);
  assign and_tmp_1 = or_612_cse & ((~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2
      | (else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[1]) | (else_7_if_div_9cyc_st_2[2])
      | (else_7_if_div_9cyc_st_2[3]));
  assign and_dcpl_3167 = ~((else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[2]));
  assign and_dcpl_3168 = and_dcpl_3167 & (~ (else_7_if_div_9cyc_st_4[3]));
  assign and_dcpl_3170 = and_1250_cse & (~ (else_7_if_div_9cyc_st_4[0]));
  assign or_tmp_23 = (max_sg1_lpi_dfm_3_st_4[15]) | (max_sg1_lpi_dfm_3_st_4[14])
      | (max_sg1_lpi_dfm_3_st_4[13]) | (max_sg1_lpi_dfm_3_st_4[0]) | (max_sg1_lpi_dfm_3_st_4[11])
      | (max_sg1_lpi_dfm_3_st_4[10]) | (max_sg1_lpi_dfm_3_st_4[9]) | (max_sg1_lpi_dfm_3_st_4[8])
      | (max_sg1_lpi_dfm_3_st_4[7]) | (max_sg1_lpi_dfm_3_st_4[6]) | (max_sg1_lpi_dfm_3_st_4[5])
      | (max_sg1_lpi_dfm_3_st_4[4]) | (max_sg1_lpi_dfm_3_st_4[3]) | (max_sg1_lpi_dfm_3_st_4[2])
      | (max_sg1_lpi_dfm_3_st_4[1]) | (max_sg1_lpi_dfm_3_st_4[12]);
  assign or_tmp_28 = (max_sg1_lpi_dfm_3_st_2[0]) | (max_sg1_lpi_dfm_3_st_2[15]) |
      (max_sg1_lpi_dfm_3_st_2[14]) | (max_sg1_lpi_dfm_3_st_2[13]) | (max_sg1_lpi_dfm_3_st_2[12])
      | (max_sg1_lpi_dfm_3_st_2[11]) | (max_sg1_lpi_dfm_3_st_2[10]) | (max_sg1_lpi_dfm_3_st_2[9])
      | (max_sg1_lpi_dfm_3_st_2[8]) | (max_sg1_lpi_dfm_3_st_2[7]) | (max_sg1_lpi_dfm_3_st_2[6])
      | (max_sg1_lpi_dfm_3_st_2[5]) | (max_sg1_lpi_dfm_3_st_2[4]) | (max_sg1_lpi_dfm_3_st_2[3])
      | (max_sg1_lpi_dfm_3_st_2[2]) | (max_sg1_lpi_dfm_3_st_2[1]);
  assign or_tmp_30 = (max_sg1_lpi_dfm_3_st_3[1]) | (max_sg1_lpi_dfm_3_st_3[15]) |
      (max_sg1_lpi_dfm_3_st_3[14]) | (max_sg1_lpi_dfm_3_st_3[13]) | (max_sg1_lpi_dfm_3_st_3[12])
      | (max_sg1_lpi_dfm_3_st_3[11]) | (max_sg1_lpi_dfm_3_st_3[10]) | (max_sg1_lpi_dfm_3_st_3[9])
      | (max_sg1_lpi_dfm_3_st_3[8]) | (max_sg1_lpi_dfm_3_st_3[7]) | (max_sg1_lpi_dfm_3_st_3[6])
      | (max_sg1_lpi_dfm_3_st_3[5]) | (max_sg1_lpi_dfm_3_st_3[4]) | (max_sg1_lpi_dfm_3_st_3[3])
      | (max_sg1_lpi_dfm_3_st_3[2]) | (max_sg1_lpi_dfm_3_st_3[0]);
  assign or_tmp_31 = (~ or_tmp_30) | (else_7_if_div_9cyc_st_3[3]) | (else_7_if_div_9cyc_st_3[2])
      | (else_7_if_div_9cyc_st_3[1]) | (else_7_if_div_9cyc_st_3[0]) | (~ main_stage_0_4)
      | if_7_equal_svs_st_3;
  assign and_dcpl_3173 = ~((else_7_if_div_9cyc_st_5[1]) | (else_7_if_div_9cyc_st_5[2]));
  assign and_dcpl_3174 = and_dcpl_3173 & (~ (else_7_if_div_9cyc_st_5[3]));
  assign and_dcpl_3176 = and_878_cse & (~ (else_7_if_div_9cyc_st_5[0]));
  assign or_tmp_33 = (max_sg1_lpi_dfm_3_st_5[0]) | (max_sg1_lpi_dfm_3_st_5[1]) |
      (max_sg1_lpi_dfm_3_st_5[2]) | (max_sg1_lpi_dfm_3_st_5[3]) | (max_sg1_lpi_dfm_3_st_5[4])
      | (max_sg1_lpi_dfm_3_st_5[5]) | (max_sg1_lpi_dfm_3_st_5[6]) | (max_sg1_lpi_dfm_3_st_5[7])
      | (max_sg1_lpi_dfm_3_st_5[8]) | (max_sg1_lpi_dfm_3_st_5[9]) | (max_sg1_lpi_dfm_3_st_5[10])
      | (max_sg1_lpi_dfm_3_st_5[11]) | (max_sg1_lpi_dfm_3_st_5[12]) | (max_sg1_lpi_dfm_3_st_5[13])
      | (max_sg1_lpi_dfm_3_st_5[14]) | (max_sg1_lpi_dfm_3_st_5[15]);
  assign or_tmp_34 = (max_sg1_lpi_dfm_3_st_4[15]) | (max_sg1_lpi_dfm_3_st_4[14])
      | (max_sg1_lpi_dfm_3_st_4[13]) | (max_sg1_lpi_dfm_3_st_4[12]) | (max_sg1_lpi_dfm_3_st_4[11])
      | (max_sg1_lpi_dfm_3_st_4[0]) | (max_sg1_lpi_dfm_3_st_4[9]) | (max_sg1_lpi_dfm_3_st_4[8])
      | (max_sg1_lpi_dfm_3_st_4[7]) | (max_sg1_lpi_dfm_3_st_4[6]) | (max_sg1_lpi_dfm_3_st_4[5])
      | (max_sg1_lpi_dfm_3_st_4[4]) | (max_sg1_lpi_dfm_3_st_4[3]) | (max_sg1_lpi_dfm_3_st_4[10])
      | (max_sg1_lpi_dfm_3_st_4[2]) | (max_sg1_lpi_dfm_3_st_4[1]);
  assign and_dcpl_3179 = ~((else_7_if_div_9cyc_st_6[1]) | (else_7_if_div_9cyc_st_6[2]));
  assign and_dcpl_3180 = and_dcpl_3179 & (~ (else_7_if_div_9cyc_st_6[3]));
  assign and_dcpl_3182 = and_506_cse & (~ (else_7_if_div_9cyc_st_6[0]));
  assign or_tmp_45 = (max_sg1_lpi_dfm_3_st_6[1]) | (max_sg1_lpi_dfm_3_st_6[0]) |
      (max_sg1_lpi_dfm_3_st_6[2]) | (max_sg1_lpi_dfm_3_st_6[3]) | (max_sg1_lpi_dfm_3_st_6[4])
      | (max_sg1_lpi_dfm_3_st_6[5]) | (max_sg1_lpi_dfm_3_st_6[6]) | (max_sg1_lpi_dfm_3_st_6[7])
      | (max_sg1_lpi_dfm_3_st_6[8]) | (max_sg1_lpi_dfm_3_st_6[9]) | (max_sg1_lpi_dfm_3_st_6[10])
      | (max_sg1_lpi_dfm_3_st_6[11]) | (max_sg1_lpi_dfm_3_st_6[12]) | (max_sg1_lpi_dfm_3_st_6[13])
      | (max_sg1_lpi_dfm_3_st_6[14]) | (max_sg1_lpi_dfm_3_st_6[15]);
  assign or_tmp_46 = (else_7_if_div_9cyc_st_5[3]) | (else_7_if_div_9cyc_st_5[2])
      | (else_7_if_div_9cyc_st_5[1]) | (else_7_if_div_9cyc_st_5[0]) | if_7_equal_svs_st_5;
  assign or_tmp_47 = (max_sg1_lpi_dfm_3_st_4[15]) | (max_sg1_lpi_dfm_3_st_4[14])
      | (max_sg1_lpi_dfm_3_st_4[13]) | (max_sg1_lpi_dfm_3_st_4[12]) | (max_sg1_lpi_dfm_3_st_4[11])
      | (max_sg1_lpi_dfm_3_st_4[10]) | (max_sg1_lpi_dfm_3_st_4[0]) | (max_sg1_lpi_dfm_3_st_4[9])
      | (max_sg1_lpi_dfm_3_st_4[8]) | (max_sg1_lpi_dfm_3_st_4[7]) | (max_sg1_lpi_dfm_3_st_4[6])
      | (max_sg1_lpi_dfm_3_st_4[5]) | (max_sg1_lpi_dfm_3_st_4[4]) | (max_sg1_lpi_dfm_3_st_4[3])
      | (max_sg1_lpi_dfm_3_st_4[2]) | (max_sg1_lpi_dfm_3_st_4[1]);
  assign and_3207_cse = ((~ or_tmp_47) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_626_cse & or_628_cse & mux_95_cse;
  assign or_tmp_58 = (max_sg1_lpi_dfm_3_st_5[15]) | (max_sg1_lpi_dfm_3_st_5[14])
      | (max_sg1_lpi_dfm_3_st_5[13]) | (max_sg1_lpi_dfm_3_st_5[12]) | (max_sg1_lpi_dfm_3_st_5[11])
      | (max_sg1_lpi_dfm_3_st_5[10]) | (max_sg1_lpi_dfm_3_st_5[9]) | (max_sg1_lpi_dfm_3_st_5[8])
      | (max_sg1_lpi_dfm_3_st_5[7]) | (max_sg1_lpi_dfm_3_st_5[6]) | (max_sg1_lpi_dfm_3_st_5[5])
      | (max_sg1_lpi_dfm_3_st_5[4]) | (max_sg1_lpi_dfm_3_st_5[3]) | (max_sg1_lpi_dfm_3_st_5[2])
      | (max_sg1_lpi_dfm_3_st_5[1]) | (max_sg1_lpi_dfm_3_st_5[0]);
  assign and_dcpl_3186 = and_dcpl_15 & (~ (else_7_if_div_9cyc_st_7[1]));
  assign and_dcpl_3188 = and_dcpl_17 & (~ (else_7_if_div_9cyc_st_7[2]));
  assign or_tmp_60 = (max_sg1_lpi_dfm_3_st_6[1]) | (max_sg1_lpi_dfm_3_st_6[2]) |
      (max_sg1_lpi_dfm_3_st_6[3]) | (max_sg1_lpi_dfm_3_st_6[4]) | (max_sg1_lpi_dfm_3_st_6[5])
      | (max_sg1_lpi_dfm_3_st_6[6]) | (max_sg1_lpi_dfm_3_st_6[7]) | (max_sg1_lpi_dfm_3_st_6[8])
      | (max_sg1_lpi_dfm_3_st_6[9]) | (max_sg1_lpi_dfm_3_st_6[10]) | (max_sg1_lpi_dfm_3_st_6[11])
      | (max_sg1_lpi_dfm_3_st_6[12]) | (max_sg1_lpi_dfm_3_st_6[13]) | (max_sg1_lpi_dfm_3_st_6[14])
      | (max_sg1_lpi_dfm_3_st_6[15]) | (max_sg1_lpi_dfm_3_st_6[0]);
  assign or_tmp_64 = (max_sg1_lpi_dfm_3_st_4[0]) | (max_sg1_lpi_dfm_3_st_4[15]) |
      (max_sg1_lpi_dfm_3_st_4[14]) | (max_sg1_lpi_dfm_3_st_4[13]) | (max_sg1_lpi_dfm_3_st_4[12])
      | (max_sg1_lpi_dfm_3_st_4[11]) | (max_sg1_lpi_dfm_3_st_4[10]) | (max_sg1_lpi_dfm_3_st_4[9])
      | (max_sg1_lpi_dfm_3_st_4[8]) | (max_sg1_lpi_dfm_3_st_4[7]) | (max_sg1_lpi_dfm_3_st_4[6])
      | (max_sg1_lpi_dfm_3_st_4[5]) | (max_sg1_lpi_dfm_3_st_4[4]) | (max_sg1_lpi_dfm_3_st_4[3])
      | (max_sg1_lpi_dfm_3_st_4[2]) | (max_sg1_lpi_dfm_3_st_4[1]);
  assign or_tmp_74 = (max_sg1_lpi_dfm_3_st_7[1]) | (max_sg1_lpi_dfm_3_st_7[3]) |
      (max_sg1_lpi_dfm_3_st_7[4]) | (max_sg1_lpi_dfm_3_st_7[5]) | (max_sg1_lpi_dfm_3_st_7[6])
      | (max_sg1_lpi_dfm_3_st_7[7]) | (max_sg1_lpi_dfm_3_st_7[8]) | (max_sg1_lpi_dfm_3_st_7[9])
      | (max_sg1_lpi_dfm_3_st_7[10]) | (max_sg1_lpi_dfm_3_st_7[11]) | (max_sg1_lpi_dfm_3_st_7[12])
      | (max_sg1_lpi_dfm_3_st_7[13]) | (max_sg1_lpi_dfm_3_st_7[14]) | (max_sg1_lpi_dfm_3_st_7[15])
      | (max_sg1_lpi_dfm_3_st_7[2]) | (max_sg1_lpi_dfm_3_st_7[0]);
  assign and_tmp_14 = or_tmp_31 & or_tmp_74;
  assign or_tmp_79 = (max_sg1_lpi_dfm_3_st_4[15]) | (max_sg1_lpi_dfm_3_st_4[14])
      | (max_sg1_lpi_dfm_3_st_4[13]) | (max_sg1_lpi_dfm_3_st_4[12]) | (max_sg1_lpi_dfm_3_st_4[11])
      | (max_sg1_lpi_dfm_3_st_4[10]) | (max_sg1_lpi_dfm_3_st_4[0]) | (max_sg1_lpi_dfm_3_st_4[8])
      | (max_sg1_lpi_dfm_3_st_4[7]) | (max_sg1_lpi_dfm_3_st_4[6]) | (max_sg1_lpi_dfm_3_st_4[5])
      | (max_sg1_lpi_dfm_3_st_4[4]) | (max_sg1_lpi_dfm_3_st_4[3]) | (max_sg1_lpi_dfm_3_st_4[2])
      | (max_sg1_lpi_dfm_3_st_4[1]) | (max_sg1_lpi_dfm_3_st_4[9]);
  assign and_tmp_22 = ((~ or_tmp_79) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_626_cse & or_628_cse & mux_95_cse;
  assign mux_102_nl = MUX_s_1_2_2({and_tmp_22 , (~(or_tmp_58 | (~ and_tmp_22)))},
      main_stage_0_6);
  assign mux_tmp_20 = MUX_s_1_2_2({(mux_102_nl) , and_tmp_22}, or_tmp_46);
  assign or_tmp_92 = (max_sg1_lpi_dfm_3_st_6[15]) | (max_sg1_lpi_dfm_3_st_6[14])
      | (max_sg1_lpi_dfm_3_st_6[13]) | (max_sg1_lpi_dfm_3_st_6[12]) | (max_sg1_lpi_dfm_3_st_6[11])
      | (max_sg1_lpi_dfm_3_st_6[10]) | (max_sg1_lpi_dfm_3_st_6[9]) | (max_sg1_lpi_dfm_3_st_6[8])
      | (max_sg1_lpi_dfm_3_st_6[7]) | (max_sg1_lpi_dfm_3_st_6[6]) | (max_sg1_lpi_dfm_3_st_6[5])
      | (max_sg1_lpi_dfm_3_st_6[4]) | (max_sg1_lpi_dfm_3_st_6[3]) | (max_sg1_lpi_dfm_3_st_6[2])
      | (max_sg1_lpi_dfm_3_st_6[1]) | (max_sg1_lpi_dfm_3_st_6[0]);
  assign mux_104_nl = MUX_s_1_2_2({mux_tmp_20 , (~(or_tmp_92 | (~ mux_tmp_20)))},
      main_stage_0_7);
  assign mux_105_cse = MUX_s_1_2_2({(mux_104_nl) , mux_tmp_20}, (else_7_if_div_9cyc_st_6[3])
      | (else_7_if_div_9cyc_st_6[2]) | (else_7_if_div_9cyc_st_6[1]) | (else_7_if_div_9cyc_st_6[0])
      | if_7_equal_svs_st_6);
  assign or_tmp_94 = (max_sg1_lpi_dfm_3_st_7[15]) | (max_sg1_lpi_dfm_3_st_7[14])
      | (max_sg1_lpi_dfm_3_st_7[13]) | (max_sg1_lpi_dfm_3_st_7[12]) | (max_sg1_lpi_dfm_3_st_7[11])
      | (max_sg1_lpi_dfm_3_st_7[10]) | (max_sg1_lpi_dfm_3_st_7[9]) | (max_sg1_lpi_dfm_3_st_7[8])
      | (max_sg1_lpi_dfm_3_st_7[7]) | (max_sg1_lpi_dfm_3_st_7[6]) | (max_sg1_lpi_dfm_3_st_7[5])
      | (max_sg1_lpi_dfm_3_st_7[4]) | (max_sg1_lpi_dfm_3_st_7[3]) | (max_sg1_lpi_dfm_3_st_7[2])
      | (max_sg1_lpi_dfm_3_st_7[1]) | (max_sg1_lpi_dfm_3_st_7[0]);
  assign and_dcpl_3238 = (~ (else_7_if_acc_tmp[1])) & (else_7_if_acc_tmp[0]);
  assign and_dcpl_3249 = (else_7_if_div_9cyc_st_2[0]) & (~ (else_7_if_div_9cyc_st_2[1]));
  assign or_tmp_184 = (else_7_if_acc_tmp[3]) | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[1])
      | (~ (else_7_if_acc_tmp[0])) | if_7_equal_tmp;
  assign or_817_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (~ (else_7_if_div_9cyc_st_1[0])) | (else_7_if_div_9cyc_st_1[1]) | (else_7_if_div_9cyc_st_1[2])
      | (else_7_if_div_9cyc_st_1[3]);
  assign and_tmp_46 = or_817_cse & or_tmp_12;
  assign and_dcpl_3258 = and_1622_cse & (else_7_if_div_9cyc_st_3[0]);
  assign and_tmp_47 = or_817_cse & ((~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2
      | (~ (else_7_if_div_9cyc_st_2[0])) | (else_7_if_div_9cyc_st_2[1]) | (else_7_if_div_9cyc_st_2[2])
      | (else_7_if_div_9cyc_st_2[3]));
  assign and_dcpl_3264 = and_1250_cse & (else_7_if_div_9cyc_st_4[0]);
  assign or_tmp_206 = (~ or_tmp_30) | (else_7_if_div_9cyc_st_3[3]) | (else_7_if_div_9cyc_st_3[2])
      | (else_7_if_div_9cyc_st_3[1]) | (~ (else_7_if_div_9cyc_st_3[0])) | (~ main_stage_0_4)
      | if_7_equal_svs_st_3;
  assign and_dcpl_3270 = and_878_cse & (else_7_if_div_9cyc_st_5[0]);
  assign and_dcpl_3276 = and_506_cse & (else_7_if_div_9cyc_st_6[0]);
  assign or_tmp_221 = (else_7_if_div_9cyc_st_5[3]) | (else_7_if_div_9cyc_st_5[2])
      | (else_7_if_div_9cyc_st_5[1]) | (~ (else_7_if_div_9cyc_st_5[0])) | if_7_equal_svs_st_5;
  assign and_3347_cse = ((~ or_tmp_47) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0])) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_831_cse & or_833_cse & mux_124_cse;
  assign and_dcpl_3280 = and_dcpl_27 & (~ (else_7_if_div_9cyc_st_7[1]));
  assign and_tmp_60 = or_tmp_206 & or_tmp_74;
  assign and_tmp_68 = ((~ or_tmp_79) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0])) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_831_cse & or_833_cse & mux_124_cse;
  assign mux_131_nl = MUX_s_1_2_2({and_tmp_68 , (~(or_tmp_58 | (~ and_tmp_68)))},
      main_stage_0_6);
  assign mux_tmp_49 = MUX_s_1_2_2({(mux_131_nl) , and_tmp_68}, or_tmp_221);
  assign mux_133_nl = MUX_s_1_2_2({mux_tmp_49 , (~(or_tmp_92 | (~ mux_tmp_49)))},
      main_stage_0_7);
  assign mux_134_cse = MUX_s_1_2_2({(mux_133_nl) , mux_tmp_49}, (else_7_if_div_9cyc_st_6[3])
      | (else_7_if_div_9cyc_st_6[2]) | (else_7_if_div_9cyc_st_6[1]) | (~ (else_7_if_div_9cyc_st_6[0]))
      | if_7_equal_svs_st_6);
  assign and_dcpl_3332 = (else_7_if_acc_tmp[1]) & (~ (else_7_if_acc_tmp[0]));
  assign and_dcpl_3337 = (~ (else_7_if_div_9cyc_st_1[2])) & (else_7_if_div_9cyc_st_1[1]);
  assign and_dcpl_3343 = (~ (else_7_if_div_9cyc_st_2[0])) & (else_7_if_div_9cyc_st_2[1]);
  assign or_tmp_359 = (else_7_if_acc_tmp[3]) | (else_7_if_acc_tmp[2]) | (~ (else_7_if_acc_tmp[1]))
      | (else_7_if_acc_tmp[0]) | if_7_equal_tmp;
  assign or_1022_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (else_7_if_div_9cyc_st_1[0]) | (~ (else_7_if_div_9cyc_st_1[1])) | (else_7_if_div_9cyc_st_1[2])
      | (else_7_if_div_9cyc_st_1[3]);
  assign and_tmp_92 = or_1022_cse & or_tmp_12;
  assign and_dcpl_3350 = (else_7_if_div_9cyc_st_3[1]) & (~ (else_7_if_div_9cyc_st_3[2]))
      & (~ (else_7_if_div_9cyc_st_3[3]));
  assign and_tmp_93 = or_1022_cse & ((~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2
      | (else_7_if_div_9cyc_st_2[0]) | (~ (else_7_if_div_9cyc_st_2[1])) | (else_7_if_div_9cyc_st_2[2])
      | (else_7_if_div_9cyc_st_2[3]));
  assign and_dcpl_3356 = (else_7_if_div_9cyc_st_4[1]) & (~ (else_7_if_div_9cyc_st_4[2]))
      & (~ (else_7_if_div_9cyc_st_4[3]));
  assign or_tmp_381 = (~ or_tmp_30) | (else_7_if_div_9cyc_st_3[3]) | (else_7_if_div_9cyc_st_3[2])
      | (~ (else_7_if_div_9cyc_st_3[1])) | (else_7_if_div_9cyc_st_3[0]) | (~ main_stage_0_4)
      | if_7_equal_svs_st_3;
  assign and_dcpl_3362 = (else_7_if_div_9cyc_st_5[1]) & (~ (else_7_if_div_9cyc_st_5[2]))
      & (~ (else_7_if_div_9cyc_st_5[3]));
  assign and_dcpl_3368 = (else_7_if_div_9cyc_st_6[1]) & (~ (else_7_if_div_9cyc_st_6[2]))
      & (~ (else_7_if_div_9cyc_st_6[3]));
  assign or_tmp_396 = (else_7_if_div_9cyc_st_5[3]) | (else_7_if_div_9cyc_st_5[2])
      | (~ (else_7_if_div_9cyc_st_5[1])) | (else_7_if_div_9cyc_st_5[0]) | if_7_equal_svs_st_5;
  assign and_3487_cse = ((~ or_tmp_47) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1036_cse & or_1038_cse & mux_153_cse;
  assign and_dcpl_3374 = and_dcpl_15 & (else_7_if_div_9cyc_st_7[1]);
  assign and_tmp_106 = or_tmp_381 & or_tmp_74;
  assign and_tmp_114 = ((~ or_tmp_79) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1036_cse & or_1038_cse & mux_153_cse;
  assign mux_160_nl = MUX_s_1_2_2({and_tmp_114 , (~(or_tmp_58 | (~ and_tmp_114)))},
      main_stage_0_6);
  assign mux_tmp_78 = MUX_s_1_2_2({(mux_160_nl) , and_tmp_114}, or_tmp_396);
  assign mux_162_nl = MUX_s_1_2_2({mux_tmp_78 , (~(or_tmp_92 | (~ mux_tmp_78)))},
      main_stage_0_7);
  assign mux_163_cse = MUX_s_1_2_2({(mux_162_nl) , mux_tmp_78}, (else_7_if_div_9cyc_st_6[3])
      | (else_7_if_div_9cyc_st_6[2]) | (~ (else_7_if_div_9cyc_st_6[1])) | (else_7_if_div_9cyc_st_6[0])
      | if_7_equal_svs_st_6);
  assign and_dcpl_3426 = (else_7_if_acc_tmp[1]) & (else_7_if_acc_tmp[0]);
  assign and_dcpl_3437 = (else_7_if_div_9cyc_st_2[0]) & (else_7_if_div_9cyc_st_2[1]);
  assign or_tmp_534 = (else_7_if_acc_tmp[3]) | (else_7_if_acc_tmp[2]) | (~ (else_7_if_acc_tmp[1]))
      | (~ (else_7_if_acc_tmp[0])) | if_7_equal_tmp;
  assign or_1227_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (~ (else_7_if_div_9cyc_st_1[0])) | (~ (else_7_if_div_9cyc_st_1[1])) | (else_7_if_div_9cyc_st_1[2])
      | (else_7_if_div_9cyc_st_1[3]);
  assign and_tmp_138 = or_1227_cse & or_tmp_12;
  assign and_tmp_139 = or_1227_cse & ((~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2
      | (~ (else_7_if_div_9cyc_st_2[0])) | (~ (else_7_if_div_9cyc_st_2[1])) | (else_7_if_div_9cyc_st_2[2])
      | (else_7_if_div_9cyc_st_2[3]));
  assign or_tmp_556 = (~ or_tmp_30) | (else_7_if_div_9cyc_st_3[3]) | (else_7_if_div_9cyc_st_3[2])
      | (~ (else_7_if_div_9cyc_st_3[1])) | (~ (else_7_if_div_9cyc_st_3[0])) | (~
      main_stage_0_4) | if_7_equal_svs_st_3;
  assign or_tmp_571 = (else_7_if_div_9cyc_st_5[3]) | (else_7_if_div_9cyc_st_5[2])
      | (~ (else_7_if_div_9cyc_st_5[1])) | (~ (else_7_if_div_9cyc_st_5[0])) | if_7_equal_svs_st_5;
  assign and_3627_cse = ((~ or_tmp_47) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (~ (else_7_if_div_9cyc_st_4[1])) | (~ (else_7_if_div_9cyc_st_4[0])) | (~
      main_stage_0_5) | if_7_equal_svs_st_4) & or_1241_cse & or_1243_cse & mux_182_cse;
  assign and_dcpl_3468 = and_dcpl_27 & (else_7_if_div_9cyc_st_7[1]);
  assign and_tmp_152 = or_tmp_556 & or_tmp_74;
  assign and_tmp_160 = ((~ or_tmp_79) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (~ (else_7_if_div_9cyc_st_4[1])) | (~ (else_7_if_div_9cyc_st_4[0])) | (~
      main_stage_0_5) | if_7_equal_svs_st_4) & or_1241_cse & or_1243_cse & mux_182_cse;
  assign mux_189_nl = MUX_s_1_2_2({and_tmp_160 , (~(or_tmp_58 | (~ and_tmp_160)))},
      main_stage_0_6);
  assign mux_tmp_107 = MUX_s_1_2_2({(mux_189_nl) , and_tmp_160}, or_tmp_571);
  assign mux_191_nl = MUX_s_1_2_2({mux_tmp_107 , (~(or_tmp_92 | (~ mux_tmp_107)))},
      main_stage_0_7);
  assign mux_192_cse = MUX_s_1_2_2({(mux_191_nl) , mux_tmp_107}, (else_7_if_div_9cyc_st_6[3])
      | (else_7_if_div_9cyc_st_6[2]) | (~ (else_7_if_div_9cyc_st_6[1])) | (~ (else_7_if_div_9cyc_st_6[0]))
      | if_7_equal_svs_st_6);
  assign and_dcpl_3522 = and_dcpl_3145 & (else_7_if_acc_tmp[2]);
  assign and_dcpl_3525 = (else_7_if_div_9cyc_st_1[2]) & (~ (else_7_if_div_9cyc_st_1[1]));
  assign or_tmp_709 = (else_7_if_acc_tmp[3]) | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[1])
      | (else_7_if_acc_tmp[0]) | if_7_equal_tmp;
  assign or_1432_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (else_7_if_div_9cyc_st_1[0]) | (else_7_if_div_9cyc_st_1[1]) | (~ (else_7_if_div_9cyc_st_1[2]))
      | (else_7_if_div_9cyc_st_1[3]);
  assign and_tmp_184 = or_1432_cse & or_tmp_12;
  assign and_dcpl_3538 = (~ (else_7_if_div_9cyc_st_3[1])) & (else_7_if_div_9cyc_st_3[2])
      & (~ (else_7_if_div_9cyc_st_3[3]));
  assign and_tmp_185 = or_1432_cse & ((~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2
      | (else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[1]) | (~ (else_7_if_div_9cyc_st_2[2]))
      | (else_7_if_div_9cyc_st_2[3]));
  assign and_dcpl_3544 = (~ (else_7_if_div_9cyc_st_4[1])) & (else_7_if_div_9cyc_st_4[2])
      & (~ (else_7_if_div_9cyc_st_4[3]));
  assign or_tmp_731 = (~ or_tmp_30) | (else_7_if_div_9cyc_st_3[3]) | (~ (else_7_if_div_9cyc_st_3[2]))
      | (else_7_if_div_9cyc_st_3[1]) | (else_7_if_div_9cyc_st_3[0]) | (~ main_stage_0_4)
      | if_7_equal_svs_st_3;
  assign and_dcpl_3550 = (~ (else_7_if_div_9cyc_st_5[1])) & (else_7_if_div_9cyc_st_5[2])
      & (~ (else_7_if_div_9cyc_st_5[3]));
  assign and_dcpl_3556 = (~ (else_7_if_div_9cyc_st_6[1])) & (else_7_if_div_9cyc_st_6[2])
      & (~ (else_7_if_div_9cyc_st_6[3]));
  assign or_tmp_746 = (else_7_if_div_9cyc_st_5[3]) | (~ (else_7_if_div_9cyc_st_5[2]))
      | (else_7_if_div_9cyc_st_5[1]) | (else_7_if_div_9cyc_st_5[0]) | if_7_equal_svs_st_5;
  assign and_3767_cse = ((~ or_tmp_47) | (else_7_if_div_9cyc_st_4[3]) | (~ (else_7_if_div_9cyc_st_4[2]))
      | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1446_cse & or_1448_cse & mux_213_cse;
  assign and_dcpl_3564 = and_dcpl_17 & (else_7_if_div_9cyc_st_7[2]);
  assign and_tmp_198 = or_tmp_731 & or_tmp_74;
  assign and_tmp_206 = ((~ or_tmp_79) | (else_7_if_div_9cyc_st_4[3]) | (~ (else_7_if_div_9cyc_st_4[2]))
      | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1446_cse & or_1448_cse & mux_213_cse;
  assign mux_220_nl = MUX_s_1_2_2({and_tmp_206 , (~(or_tmp_58 | (~ and_tmp_206)))},
      main_stage_0_6);
  assign mux_tmp_138 = MUX_s_1_2_2({(mux_220_nl) , and_tmp_206}, or_tmp_746);
  assign mux_222_nl = MUX_s_1_2_2({mux_tmp_138 , (~(or_tmp_92 | (~ mux_tmp_138)))},
      main_stage_0_7);
  assign mux_223_cse = MUX_s_1_2_2({(mux_222_nl) , mux_tmp_138}, (else_7_if_div_9cyc_st_6[3])
      | (~ (else_7_if_div_9cyc_st_6[2])) | (else_7_if_div_9cyc_st_6[1]) | (else_7_if_div_9cyc_st_6[0])
      | if_7_equal_svs_st_6);
  assign or_tmp_884 = (else_7_if_acc_tmp[3]) | (~ (else_7_if_acc_tmp[2])) | (else_7_if_acc_tmp[1])
      | (~ (else_7_if_acc_tmp[0])) | if_7_equal_tmp;
  assign or_1637_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (~ (else_7_if_div_9cyc_st_1[0])) | (else_7_if_div_9cyc_st_1[1]) | (~ (else_7_if_div_9cyc_st_1[2]))
      | (else_7_if_div_9cyc_st_1[3]);
  assign and_tmp_230 = or_1637_cse & or_tmp_12;
  assign and_tmp_231 = or_1637_cse & ((~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2
      | (~ (else_7_if_div_9cyc_st_2[0])) | (else_7_if_div_9cyc_st_2[1]) | (~ (else_7_if_div_9cyc_st_2[2]))
      | (else_7_if_div_9cyc_st_2[3]));
  assign or_tmp_906 = (~ or_tmp_30) | (else_7_if_div_9cyc_st_3[3]) | (~ (else_7_if_div_9cyc_st_3[2]))
      | (else_7_if_div_9cyc_st_3[1]) | (~ (else_7_if_div_9cyc_st_3[0])) | (~ main_stage_0_4)
      | if_7_equal_svs_st_3;
  assign or_tmp_921 = (else_7_if_div_9cyc_st_5[3]) | (~ (else_7_if_div_9cyc_st_5[2]))
      | (else_7_if_div_9cyc_st_5[1]) | (~ (else_7_if_div_9cyc_st_5[0])) | if_7_equal_svs_st_5;
  assign and_3907_cse = ((~ or_tmp_47) | (else_7_if_div_9cyc_st_4[3]) | (~ (else_7_if_div_9cyc_st_4[2]))
      | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0])) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1651_cse & or_1653_cse & mux_242_cse;
  assign and_tmp_244 = or_tmp_906 & or_tmp_74;
  assign and_tmp_252 = ((~ or_tmp_79) | (else_7_if_div_9cyc_st_4[3]) | (~ (else_7_if_div_9cyc_st_4[2]))
      | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0])) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1651_cse & or_1653_cse & mux_242_cse;
  assign mux_249_nl = MUX_s_1_2_2({and_tmp_252 , (~(or_tmp_58 | (~ and_tmp_252)))},
      main_stage_0_6);
  assign mux_tmp_167 = MUX_s_1_2_2({(mux_249_nl) , and_tmp_252}, or_tmp_921);
  assign mux_251_nl = MUX_s_1_2_2({mux_tmp_167 , (~(or_tmp_92 | (~ mux_tmp_167)))},
      main_stage_0_7);
  assign mux_252_cse = MUX_s_1_2_2({(mux_251_nl) , mux_tmp_167}, (else_7_if_div_9cyc_st_6[3])
      | (~ (else_7_if_div_9cyc_st_6[2])) | (else_7_if_div_9cyc_st_6[1]) | (~ (else_7_if_div_9cyc_st_6[0]))
      | if_7_equal_svs_st_6);
  assign and_dcpl_3713 = (else_7_if_div_9cyc_st_1[2]) & (else_7_if_div_9cyc_st_1[1]);
  assign or_tmp_1059 = (else_7_if_acc_tmp[3]) | (~ (else_7_if_acc_tmp[2])) | (~ (else_7_if_acc_tmp[1]))
      | (else_7_if_acc_tmp[0]) | if_7_equal_tmp;
  assign or_1842_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (else_7_if_div_9cyc_st_1[0]) | (~ (else_7_if_div_9cyc_st_1[1])) | (~ (else_7_if_div_9cyc_st_1[2]))
      | (else_7_if_div_9cyc_st_1[3]);
  assign and_tmp_276 = or_1842_cse & or_tmp_12;
  assign and_dcpl_3726 = (else_7_if_div_9cyc_st_3[1]) & (else_7_if_div_9cyc_st_3[2])
      & (~ (else_7_if_div_9cyc_st_3[3]));
  assign and_tmp_277 = or_1842_cse & ((~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2
      | (else_7_if_div_9cyc_st_2[0]) | (~ (else_7_if_div_9cyc_st_2[1])) | (~ (else_7_if_div_9cyc_st_2[2]))
      | (else_7_if_div_9cyc_st_2[3]));
  assign and_dcpl_3732 = (else_7_if_div_9cyc_st_4[1]) & (else_7_if_div_9cyc_st_4[2])
      & (~ (else_7_if_div_9cyc_st_4[3]));
  assign or_tmp_1081 = (~ or_tmp_30) | (else_7_if_div_9cyc_st_3[3]) | (~ (else_7_if_div_9cyc_st_3[2]))
      | (~ (else_7_if_div_9cyc_st_3[1])) | (else_7_if_div_9cyc_st_3[0]) | (~ main_stage_0_4)
      | if_7_equal_svs_st_3;
  assign and_dcpl_3738 = (else_7_if_div_9cyc_st_5[1]) & (else_7_if_div_9cyc_st_5[2])
      & (~ (else_7_if_div_9cyc_st_5[3]));
  assign and_dcpl_3744 = (else_7_if_div_9cyc_st_6[1]) & (else_7_if_div_9cyc_st_6[2])
      & (~ (else_7_if_div_9cyc_st_6[3]));
  assign or_tmp_1096 = (else_7_if_div_9cyc_st_5[3]) | (~ (else_7_if_div_9cyc_st_5[2]))
      | (~ (else_7_if_div_9cyc_st_5[1])) | (else_7_if_div_9cyc_st_5[0]) | if_7_equal_svs_st_5;
  assign and_4047_cse = ((~ or_tmp_47) | (else_7_if_div_9cyc_st_4[3]) | (~ (else_7_if_div_9cyc_st_4[2]))
      | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1856_cse & or_1858_cse & mux_271_cse;
  assign and_tmp_290 = or_tmp_1081 & or_tmp_74;
  assign and_tmp_298 = ((~ or_tmp_79) | (else_7_if_div_9cyc_st_4[3]) | (~ (else_7_if_div_9cyc_st_4[2]))
      | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1856_cse & or_1858_cse & mux_271_cse;
  assign mux_278_nl = MUX_s_1_2_2({and_tmp_298 , (~(or_tmp_58 | (~ and_tmp_298)))},
      main_stage_0_6);
  assign mux_tmp_196 = MUX_s_1_2_2({(mux_278_nl) , and_tmp_298}, or_tmp_1096);
  assign mux_280_nl = MUX_s_1_2_2({mux_tmp_196 , (~(or_tmp_92 | (~ mux_tmp_196)))},
      main_stage_0_7);
  assign mux_281_cse = MUX_s_1_2_2({(mux_280_nl) , mux_tmp_196}, (else_7_if_div_9cyc_st_6[3])
      | (~ (else_7_if_div_9cyc_st_6[2])) | (~ (else_7_if_div_9cyc_st_6[1])) | (else_7_if_div_9cyc_st_6[0])
      | if_7_equal_svs_st_6);
  assign or_tmp_1234 = (else_7_if_acc_tmp[3]) | (~ (else_7_if_acc_tmp[2])) | (~ (else_7_if_acc_tmp[1]))
      | (~ (else_7_if_acc_tmp[0])) | if_7_equal_tmp;
  assign nand_cse = ~(or_tmp_10 & main_stage_0_2 & (~ if_7_equal_svs_st_1) & (else_7_if_div_9cyc_st_1[0])
      & (else_7_if_div_9cyc_st_1[1]) & (else_7_if_div_9cyc_st_1[2]) & (~ (else_7_if_div_9cyc_st_1[3])));
  assign and_tmp_322 = nand_cse & or_tmp_12;
  assign and_tmp_323 = nand_cse & (~(or_tmp_12 & main_stage_0_3 & (~ if_7_equal_svs_st_2)
      & (else_7_if_div_9cyc_st_2[0]) & (else_7_if_div_9cyc_st_2[1]) & (else_7_if_div_9cyc_st_2[2])
      & (~ (else_7_if_div_9cyc_st_2[3]))));
  assign or_tmp_1256 = ~(or_tmp_30 & (~ (else_7_if_div_9cyc_st_3[3])) & (else_7_if_div_9cyc_st_3[2])
      & (else_7_if_div_9cyc_st_3[1]) & (else_7_if_div_9cyc_st_3[0]) & main_stage_0_4
      & (~ if_7_equal_svs_st_3));
  assign or_tmp_1271 = (else_7_if_div_9cyc_st_5[3]) | (~ (else_7_if_div_9cyc_st_5[2]))
      | (~ (else_7_if_div_9cyc_st_5[1])) | (~ (else_7_if_div_9cyc_st_5[0])) | if_7_equal_svs_st_5;
  assign mux_302_cse = MUX_s_1_2_2({(~(main_stage_0_3 | (~ or_tmp_1256))) , or_tmp_1256},
      or_2065_cse);
  assign and_4187_cse = (~(or_tmp_47 & (~ (else_7_if_div_9cyc_st_4[3])) & (else_7_if_div_9cyc_st_4[2])
      & (else_7_if_div_9cyc_st_4[1]) & (else_7_if_div_9cyc_st_4[0]) & main_stage_0_5
      & (~ if_7_equal_svs_st_4))) & or_2061_cse & nand_33_cse & mux_302_cse;
  assign and_4195_cse = or_tmp_1256 & or_tmp_74;
  assign and_tmp_344 = (~(or_tmp_79 & (~ (else_7_if_div_9cyc_st_4[3])) & (else_7_if_div_9cyc_st_4[2])
      & (else_7_if_div_9cyc_st_4[1]) & (else_7_if_div_9cyc_st_4[0]) & main_stage_0_5
      & (~ if_7_equal_svs_st_4))) & or_2061_cse & nand_33_cse & mux_302_cse;
  assign mux_307_nl = MUX_s_1_2_2({and_tmp_344 , (~(or_tmp_58 | (~ and_tmp_344)))},
      main_stage_0_6);
  assign mux_tmp_225 = MUX_s_1_2_2({(mux_307_nl) , and_tmp_344}, or_tmp_1271);
  assign mux_309_nl = MUX_s_1_2_2({mux_tmp_225 , (~(or_tmp_92 | (~ mux_tmp_225)))},
      main_stage_0_7);
  assign mux_310_cse = MUX_s_1_2_2({(mux_309_nl) , mux_tmp_225}, (else_7_if_div_9cyc_st_6[3])
      | (~ (else_7_if_div_9cyc_st_6[2])) | (~ (else_7_if_div_9cyc_st_6[1])) | (~
      (else_7_if_div_9cyc_st_6[0])) | if_7_equal_svs_st_6);
  assign or_tmp_1409 = (~ (else_7_if_acc_tmp[3])) | (else_7_if_acc_tmp[2]) | (else_7_if_acc_tmp[1])
      | (else_7_if_acc_tmp[0]) | if_7_equal_tmp;
  assign or_2252_cse = (~ or_tmp_10) | (~ main_stage_0_2) | if_7_equal_svs_st_1 |
      (else_7_if_div_9cyc_st_1[0]) | (else_7_if_div_9cyc_st_1[1]) | (else_7_if_div_9cyc_st_1[2]);
  assign mux_tmp_246 = MUX_s_1_2_2({(~((else_7_if_div_9cyc_st_1[3]) | (~ or_tmp_12)))
      , or_tmp_12}, or_2252_cse);
  assign or_tmp_1422 = (~ or_tmp_12) | (~ main_stage_0_3) | if_7_equal_svs_st_2 |
      (else_7_if_div_9cyc_st_2[0]) | (else_7_if_div_9cyc_st_2[1]) | (else_7_if_div_9cyc_st_2[2])
      | (~ (else_7_if_div_9cyc_st_2[3]));
  assign mux_tmp_248 = MUX_s_1_2_2({(~((else_7_if_div_9cyc_st_1[3]) | (~ or_tmp_1422)))
      , or_tmp_1422}, or_2252_cse);
  assign or_tmp_1434 = (~ or_tmp_30) | (~ (else_7_if_div_9cyc_st_3[3])) | (else_7_if_div_9cyc_st_3[2])
      | (else_7_if_div_9cyc_st_3[1]) | (else_7_if_div_9cyc_st_3[0]) | (~ main_stage_0_4)
      | if_7_equal_svs_st_3;
  assign or_tmp_1449 = (~ (else_7_if_div_9cyc_st_5[3])) | (else_7_if_div_9cyc_st_5[2])
      | (else_7_if_div_9cyc_st_5[1]) | (else_7_if_div_9cyc_st_5[0]) | if_7_equal_svs_st_5;
  assign and_4325_cse = ((~ or_tmp_47) | (~ (else_7_if_div_9cyc_st_4[3])) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_2269_cse & or_2271_cse & mux_333_cse;
  assign and_tmp_380 = or_tmp_1434 & or_tmp_74;
  assign and_tmp_388 = ((~ or_tmp_79) | (~ (else_7_if_div_9cyc_st_4[3])) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_2269_cse & or_2271_cse & mux_333_cse;
  assign mux_340_nl = MUX_s_1_2_2({and_tmp_388 , (~(or_tmp_58 | (~ and_tmp_388)))},
      main_stage_0_6);
  assign mux_tmp_258 = MUX_s_1_2_2({(mux_340_nl) , and_tmp_388}, or_tmp_1449);
  assign mux_342_nl = MUX_s_1_2_2({mux_tmp_258 , (~(or_tmp_92 | (~ mux_tmp_258)))},
      main_stage_0_7);
  assign mux_343_cse = MUX_s_1_2_2({(mux_342_nl) , mux_tmp_258}, (~ (else_7_if_div_9cyc_st_6[3]))
      | (else_7_if_div_9cyc_st_6[2]) | (else_7_if_div_9cyc_st_6[1]) | (else_7_if_div_9cyc_st_6[0])
      | if_7_equal_svs_st_6);
  assign and_dcpl_3990 = ~((else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[0]));
  assign and_dcpl_3991 = and_dcpl_3990 & (~ (else_7_if_1_acc_tmp[2]));
  assign and_dcpl_3992 = (~ if_7_equal_tmp) & else_7_equal_tmp;
  assign and_dcpl_3993 = and_dcpl_3992 & (~ (else_7_if_1_acc_tmp[1]));
  assign and_dcpl_3996 = and_dcpl_2356 & (~ (else_7_if_1_div_9cyc[0]));
  assign and_dcpl_3997 = main_stage_0_2 & else_7_equal_svs_st_1;
  assign and_dcpl_3998 = and_dcpl_3997 & (~ (else_7_if_1_div_9cyc[2]));
  assign or_dcpl_854 = (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[0]);
  assign or_dcpl_855 = or_dcpl_854 | (else_7_if_1_acc_tmp[2]);
  assign or_dcpl_856 = if_7_equal_tmp | (~ else_7_equal_tmp);
  assign or_dcpl_857 = or_dcpl_856 | (else_7_if_1_acc_tmp[1]);
  assign and_dcpl_4003 = and_dcpl_1984 & (~ (else_7_if_1_div_9cyc_st_2[0]));
  assign and_dcpl_4006 = and_1994_cse & else_7_equal_svs_st_2 & (~ (else_7_if_1_div_9cyc_st_2[2]));
  assign and_dcpl_4010 = and_dcpl_1612 & (~ (else_7_if_1_div_9cyc_st_3[2]));
  assign and_dcpl_4013 = and_1622_cse & else_7_equal_svs_st_3 & (~ (else_7_if_1_div_9cyc_st_3[0]));
  assign or_tmp_1591 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_9cyc_st_2[0]) | (else_7_if_1_div_9cyc_st_2[1]) | (else_7_if_1_div_9cyc_st_2[2])
      | (else_7_if_1_div_9cyc_st_2[3]);
  assign or_tmp_1592 = (else_7_if_1_div_9cyc[0]) | (else_7_if_1_div_9cyc[1]) | (else_7_if_1_div_9cyc[2])
      | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2) | if_7_equal_svs_st_1;
  assign or_tmp_1593 = (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[2]) | (else_7_if_1_acc_tmp[1])
      | (else_7_if_1_acc_tmp[0]) | (~ else_7_equal_tmp) | if_7_equal_tmp;
  assign and_dcpl_4017 = and_dcpl_1240 & (~ (else_7_if_1_div_9cyc_st_4[1]));
  assign and_dcpl_4020 = and_1250_cse & else_7_equal_svs_st_4 & (~ (else_7_if_1_div_9cyc_st_4[2]));
  assign or_tmp_1595 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (else_7_if_1_div_9cyc_st_3[0]) | (else_7_if_1_div_9cyc_st_3[1]) | (else_7_if_1_div_9cyc_st_3[2])
      | (else_7_if_1_div_9cyc_st_3[3]);
  assign and_dcpl_4024 = and_dcpl_868 & (~ (else_7_if_1_div_9cyc_st_5[0]));
  assign and_dcpl_4027 = and_878_cse & else_7_equal_svs_st_5 & (~ (else_7_if_1_div_9cyc_st_5[3]));
  assign or_tmp_1600 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (else_7_if_1_div_9cyc_st_4[0]) | (else_7_if_1_div_9cyc_st_4[1]) | (else_7_if_1_div_9cyc_st_4[2])
      | (else_7_if_1_div_9cyc_st_4[3]);
  assign and_dcpl_4031 = and_dcpl_496 & (~ (else_7_if_1_div_9cyc_st_6[1]));
  assign and_dcpl_4034 = and_506_cse & else_7_equal_svs_st_6 & (~ (else_7_if_1_div_9cyc_st_6[2]));
  assign or_tmp_1606 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (else_7_if_1_div_9cyc_st_5[0]) | (else_7_if_1_div_9cyc_st_5[1]) | (else_7_if_1_div_9cyc_st_5[2])
      | (else_7_if_1_div_9cyc_st_5[3]);
  assign and_dcpl_4038 = and_dcpl_124 & (~ (else_7_if_1_div_9cyc_st_7[1]));
  assign and_dcpl_4041 = and_dcpl_17 & else_7_equal_svs_st_7 & (~ (else_7_if_1_div_9cyc_st_7[2]));
  assign or_tmp_1613 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (else_7_if_1_div_9cyc_st_6[0]) | (else_7_if_1_div_9cyc_st_6[1]) | (else_7_if_1_div_9cyc_st_6[2])
      | (else_7_if_1_div_9cyc_st_6[3]);
  assign and_tmp_421 = or_tmp_1593 & or_tmp_1591;
  assign and_dcpl_4098 = (~ (else_7_if_1_acc_tmp[3])) & (else_7_if_1_acc_tmp[0]);
  assign and_dcpl_4099 = and_dcpl_4098 & (~ (else_7_if_1_acc_tmp[2]));
  assign and_dcpl_4104 = and_dcpl_2356 & (else_7_if_1_div_9cyc[0]);
  assign or_dcpl_864 = (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[0]));
  assign or_dcpl_865 = or_dcpl_864 | (else_7_if_1_acc_tmp[2]);
  assign and_dcpl_4111 = and_dcpl_1984 & (else_7_if_1_div_9cyc_st_2[0]);
  assign and_dcpl_4121 = and_1622_cse & else_7_equal_svs_st_3 & (else_7_if_1_div_9cyc_st_3[0]);
  assign or_tmp_1671 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (~ (else_7_if_1_div_9cyc_st_2[0])) | (else_7_if_1_div_9cyc_st_2[1]) | (else_7_if_1_div_9cyc_st_2[2])
      | (else_7_if_1_div_9cyc_st_2[3]);
  assign or_tmp_1672 = (~ (else_7_if_1_div_9cyc[0])) | (else_7_if_1_div_9cyc[1])
      | (else_7_if_1_div_9cyc[2]) | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_tmp_1673 = (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[2]) | (else_7_if_1_acc_tmp[1])
      | (~ (else_7_if_1_acc_tmp[0])) | (~ else_7_equal_tmp) | if_7_equal_tmp;
  assign and_dcpl_4125 = and_dcpl_1252 & (~ (else_7_if_1_div_9cyc_st_4[1]));
  assign or_tmp_1675 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (~ (else_7_if_1_div_9cyc_st_3[0])) | (else_7_if_1_div_9cyc_st_3[1]) | (else_7_if_1_div_9cyc_st_3[2])
      | (else_7_if_1_div_9cyc_st_3[3]);
  assign or_tmp_1680 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (~ (else_7_if_1_div_9cyc_st_4[0])) | (else_7_if_1_div_9cyc_st_4[1]) | (else_7_if_1_div_9cyc_st_4[2])
      | (else_7_if_1_div_9cyc_st_4[3]);
  assign and_dcpl_4139 = and_dcpl_508 & (~ (else_7_if_1_div_9cyc_st_6[1]));
  assign or_tmp_1686 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (~ (else_7_if_1_div_9cyc_st_5[0])) | (else_7_if_1_div_9cyc_st_5[1]) | (else_7_if_1_div_9cyc_st_5[2])
      | (else_7_if_1_div_9cyc_st_5[3]);
  assign and_dcpl_4146 = and_dcpl_136 & (~ (else_7_if_1_div_9cyc_st_7[1]));
  assign or_tmp_1693 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (~ (else_7_if_1_div_9cyc_st_6[0])) | (else_7_if_1_div_9cyc_st_6[1]) | (else_7_if_1_div_9cyc_st_6[2])
      | (else_7_if_1_div_9cyc_st_6[3]);
  assign and_tmp_464 = or_tmp_1673 & or_tmp_1671;
  assign and_dcpl_4209 = and_dcpl_3992 & (else_7_if_1_acc_tmp[1]);
  assign and_dcpl_4212 = and_dcpl_2380 & (~ (else_7_if_1_div_9cyc[0]));
  assign or_dcpl_877 = or_dcpl_856 | (~ (else_7_if_1_acc_tmp[1]));
  assign and_dcpl_4219 = and_dcpl_2008 & (~ (else_7_if_1_div_9cyc_st_2[0]));
  assign and_dcpl_4226 = and_dcpl_1636 & (~ (else_7_if_1_div_9cyc_st_3[2]));
  assign or_tmp_1751 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_9cyc_st_2[0]) | (~ (else_7_if_1_div_9cyc_st_2[1])) | (else_7_if_1_div_9cyc_st_2[2])
      | (else_7_if_1_div_9cyc_st_2[3]);
  assign or_tmp_1752 = (else_7_if_1_div_9cyc[0]) | (~ (else_7_if_1_div_9cyc[1]))
      | (else_7_if_1_div_9cyc[2]) | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_tmp_1753 = (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[2]) | (~ (else_7_if_1_acc_tmp[1]))
      | (else_7_if_1_acc_tmp[0]) | (~ else_7_equal_tmp) | if_7_equal_tmp;
  assign and_dcpl_4233 = and_dcpl_1240 & (else_7_if_1_div_9cyc_st_4[1]);
  assign or_tmp_1755 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (else_7_if_1_div_9cyc_st_3[0]) | (~ (else_7_if_1_div_9cyc_st_3[1])) | (else_7_if_1_div_9cyc_st_3[2])
      | (else_7_if_1_div_9cyc_st_3[3]);
  assign or_tmp_1760 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (else_7_if_1_div_9cyc_st_4[0]) | (~ (else_7_if_1_div_9cyc_st_4[1])) | (else_7_if_1_div_9cyc_st_4[2])
      | (else_7_if_1_div_9cyc_st_4[3]);
  assign and_dcpl_4247 = and_dcpl_496 & (else_7_if_1_div_9cyc_st_6[1]);
  assign or_tmp_1766 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (else_7_if_1_div_9cyc_st_5[0]) | (~ (else_7_if_1_div_9cyc_st_5[1])) | (else_7_if_1_div_9cyc_st_5[2])
      | (else_7_if_1_div_9cyc_st_5[3]);
  assign and_dcpl_4254 = and_dcpl_124 & (else_7_if_1_div_9cyc_st_7[1]);
  assign or_tmp_1773 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (else_7_if_1_div_9cyc_st_6[0]) | (~ (else_7_if_1_div_9cyc_st_6[1])) | (else_7_if_1_div_9cyc_st_6[2])
      | (else_7_if_1_div_9cyc_st_6[3]);
  assign and_tmp_507 = or_tmp_1753 & or_tmp_1751;
  assign and_dcpl_4320 = and_dcpl_2380 & (else_7_if_1_div_9cyc[0]);
  assign and_dcpl_4327 = and_dcpl_2008 & (else_7_if_1_div_9cyc_st_2[0]);
  assign or_tmp_1831 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (~ (else_7_if_1_div_9cyc_st_2[0])) | (~ (else_7_if_1_div_9cyc_st_2[1])) |
      (else_7_if_1_div_9cyc_st_2[2]) | (else_7_if_1_div_9cyc_st_2[3]);
  assign or_tmp_1832 = (~ (else_7_if_1_div_9cyc[0])) | (~ (else_7_if_1_div_9cyc[1]))
      | (else_7_if_1_div_9cyc[2]) | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_tmp_1833 = (else_7_if_1_acc_tmp[3]) | (else_7_if_1_acc_tmp[2]) | (~ (else_7_if_1_acc_tmp[1]))
      | (~ (else_7_if_1_acc_tmp[0])) | (~ else_7_equal_tmp) | if_7_equal_tmp;
  assign and_dcpl_4341 = and_dcpl_1252 & (else_7_if_1_div_9cyc_st_4[1]);
  assign or_tmp_1835 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (~ (else_7_if_1_div_9cyc_st_3[0])) | (~ (else_7_if_1_div_9cyc_st_3[1])) |
      (else_7_if_1_div_9cyc_st_3[2]) | (else_7_if_1_div_9cyc_st_3[3]);
  assign or_tmp_1840 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (~ (else_7_if_1_div_9cyc_st_4[0])) | (~ (else_7_if_1_div_9cyc_st_4[1])) |
      (else_7_if_1_div_9cyc_st_4[2]) | (else_7_if_1_div_9cyc_st_4[3]);
  assign and_dcpl_4355 = and_dcpl_508 & (else_7_if_1_div_9cyc_st_6[1]);
  assign or_tmp_1846 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (~ (else_7_if_1_div_9cyc_st_5[0])) | (~ (else_7_if_1_div_9cyc_st_5[1])) |
      (else_7_if_1_div_9cyc_st_5[2]) | (else_7_if_1_div_9cyc_st_5[3]);
  assign and_dcpl_4362 = and_dcpl_136 & (else_7_if_1_div_9cyc_st_7[1]);
  assign or_tmp_1853 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (~ (else_7_if_1_div_9cyc_st_6[0])) | (~ (else_7_if_1_div_9cyc_st_6[1])) |
      (else_7_if_1_div_9cyc_st_6[2]) | (else_7_if_1_div_9cyc_st_6[3]);
  assign and_tmp_550 = or_tmp_1833 & or_tmp_1831;
  assign and_dcpl_4423 = and_dcpl_3990 & (else_7_if_1_acc_tmp[2]);
  assign and_dcpl_4430 = and_dcpl_3997 & (else_7_if_1_div_9cyc[2]);
  assign or_dcpl_895 = or_dcpl_854 | (~ (else_7_if_1_acc_tmp[2]));
  assign and_dcpl_4438 = and_1994_cse & else_7_equal_svs_st_2 & (else_7_if_1_div_9cyc_st_2[2]);
  assign and_dcpl_4442 = and_dcpl_1612 & (else_7_if_1_div_9cyc_st_3[2]);
  assign or_tmp_1911 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_9cyc_st_2[0]) | (else_7_if_1_div_9cyc_st_2[1]) | (~ (else_7_if_1_div_9cyc_st_2[2]))
      | (else_7_if_1_div_9cyc_st_2[3]);
  assign or_tmp_1912 = (else_7_if_1_div_9cyc[0]) | (else_7_if_1_div_9cyc[1]) | (~
      (else_7_if_1_div_9cyc[2])) | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_tmp_1913 = (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[2])) |
      (else_7_if_1_acc_tmp[1]) | (else_7_if_1_acc_tmp[0]) | (~ else_7_equal_tmp)
      | if_7_equal_tmp;
  assign and_dcpl_4452 = and_1250_cse & else_7_equal_svs_st_4 & (else_7_if_1_div_9cyc_st_4[2]);
  assign or_tmp_1915 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (else_7_if_1_div_9cyc_st_3[0]) | (else_7_if_1_div_9cyc_st_3[1]) | (~ (else_7_if_1_div_9cyc_st_3[2]))
      | (else_7_if_1_div_9cyc_st_3[3]);
  assign or_tmp_1920 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (else_7_if_1_div_9cyc_st_4[0]) | (else_7_if_1_div_9cyc_st_4[1]) | (~ (else_7_if_1_div_9cyc_st_4[2]))
      | (else_7_if_1_div_9cyc_st_4[3]);
  assign and_dcpl_4466 = and_506_cse & else_7_equal_svs_st_6 & (else_7_if_1_div_9cyc_st_6[2]);
  assign or_tmp_1926 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (else_7_if_1_div_9cyc_st_5[0]) | (else_7_if_1_div_9cyc_st_5[1]) | (~ (else_7_if_1_div_9cyc_st_5[2]))
      | (else_7_if_1_div_9cyc_st_5[3]);
  assign and_dcpl_4473 = and_dcpl_17 & else_7_equal_svs_st_7 & (else_7_if_1_div_9cyc_st_7[2]);
  assign or_tmp_1933 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (else_7_if_1_div_9cyc_st_6[0]) | (else_7_if_1_div_9cyc_st_6[1]) | (~ (else_7_if_1_div_9cyc_st_6[2]))
      | (else_7_if_1_div_9cyc_st_6[3]);
  assign and_tmp_593 = or_tmp_1913 & or_tmp_1911;
  assign and_dcpl_4531 = and_dcpl_4098 & (else_7_if_1_acc_tmp[2]);
  assign or_dcpl_905 = or_dcpl_864 | (~ (else_7_if_1_acc_tmp[2]));
  assign or_tmp_1991 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (~ (else_7_if_1_div_9cyc_st_2[0])) | (else_7_if_1_div_9cyc_st_2[1]) | (~
      (else_7_if_1_div_9cyc_st_2[2])) | (else_7_if_1_div_9cyc_st_2[3]);
  assign or_tmp_1992 = (~ (else_7_if_1_div_9cyc[0])) | (else_7_if_1_div_9cyc[1])
      | (~ (else_7_if_1_div_9cyc[2])) | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_tmp_1993 = (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[2])) |
      (else_7_if_1_acc_tmp[1]) | (~ (else_7_if_1_acc_tmp[0])) | (~ else_7_equal_tmp)
      | if_7_equal_tmp;
  assign or_tmp_1995 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (~ (else_7_if_1_div_9cyc_st_3[0])) | (else_7_if_1_div_9cyc_st_3[1]) | (~
      (else_7_if_1_div_9cyc_st_3[2])) | (else_7_if_1_div_9cyc_st_3[3]);
  assign or_tmp_2000 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (~ (else_7_if_1_div_9cyc_st_4[0])) | (else_7_if_1_div_9cyc_st_4[1]) | (~
      (else_7_if_1_div_9cyc_st_4[2])) | (else_7_if_1_div_9cyc_st_4[3]);
  assign or_tmp_2006 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (~ (else_7_if_1_div_9cyc_st_5[0])) | (else_7_if_1_div_9cyc_st_5[1]) | (~
      (else_7_if_1_div_9cyc_st_5[2])) | (else_7_if_1_div_9cyc_st_5[3]);
  assign or_tmp_2013 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (~ (else_7_if_1_div_9cyc_st_6[0])) | (else_7_if_1_div_9cyc_st_6[1]) | (~
      (else_7_if_1_div_9cyc_st_6[2])) | (else_7_if_1_div_9cyc_st_6[3]);
  assign and_tmp_636 = or_tmp_1993 & or_tmp_1991;
  assign and_dcpl_4658 = and_dcpl_1636 & (else_7_if_1_div_9cyc_st_3[2]);
  assign or_tmp_2071 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_9cyc_st_2[0]) | (~ (else_7_if_1_div_9cyc_st_2[1])) | (~
      (else_7_if_1_div_9cyc_st_2[2])) | (else_7_if_1_div_9cyc_st_2[3]);
  assign or_tmp_2072 = (else_7_if_1_div_9cyc[0]) | (~ (else_7_if_1_div_9cyc[1]))
      | (~ (else_7_if_1_div_9cyc[2])) | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_tmp_2073 = (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[2])) |
      (~ (else_7_if_1_acc_tmp[1])) | (else_7_if_1_acc_tmp[0]) | (~ else_7_equal_tmp)
      | if_7_equal_tmp;
  assign or_tmp_2075 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (else_7_if_1_div_9cyc_st_3[0]) | (~ (else_7_if_1_div_9cyc_st_3[1])) | (~
      (else_7_if_1_div_9cyc_st_3[2])) | (else_7_if_1_div_9cyc_st_3[3]);
  assign or_tmp_2080 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (else_7_if_1_div_9cyc_st_4[0]) | (~ (else_7_if_1_div_9cyc_st_4[1])) | (~
      (else_7_if_1_div_9cyc_st_4[2])) | (else_7_if_1_div_9cyc_st_4[3]);
  assign or_tmp_2086 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (else_7_if_1_div_9cyc_st_5[0]) | (~ (else_7_if_1_div_9cyc_st_5[1])) | (~
      (else_7_if_1_div_9cyc_st_5[2])) | (else_7_if_1_div_9cyc_st_5[3]);
  assign or_tmp_2093 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (else_7_if_1_div_9cyc_st_6[0]) | (~ (else_7_if_1_div_9cyc_st_6[1])) | (~
      (else_7_if_1_div_9cyc_st_6[2])) | (else_7_if_1_div_9cyc_st_6[3]);
  assign and_tmp_679 = or_tmp_2073 & or_tmp_2071;
  assign or_tmp_2151 = ~(main_stage_0_3 & (~ if_7_equal_svs_st_2) & else_7_equal_svs_st_2
      & (else_7_if_1_div_9cyc_st_2[0]) & (else_7_if_1_div_9cyc_st_2[1]) & (else_7_if_1_div_9cyc_st_2[2])
      & (~ (else_7_if_1_div_9cyc_st_2[3])));
  assign or_tmp_2152 = (~ (else_7_if_1_div_9cyc[0])) | (~ (else_7_if_1_div_9cyc[1]))
      | (~ (else_7_if_1_div_9cyc[2])) | (else_7_if_1_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1;
  assign or_tmp_2153 = (else_7_if_1_acc_tmp[3]) | (~ (else_7_if_1_acc_tmp[2])) |
      (~ (else_7_if_1_acc_tmp[1])) | (~ (else_7_if_1_acc_tmp[0])) | (~ else_7_equal_tmp)
      | if_7_equal_tmp;
  assign or_tmp_2155 = ~(main_stage_0_4 & (~ if_7_equal_svs_st_3) & else_7_equal_svs_st_3
      & (else_7_if_1_div_9cyc_st_3[0]) & (else_7_if_1_div_9cyc_st_3[1]) & (else_7_if_1_div_9cyc_st_3[2])
      & (~ (else_7_if_1_div_9cyc_st_3[3])));
  assign or_tmp_2160 = ~(main_stage_0_5 & (~ if_7_equal_svs_st_4) & else_7_equal_svs_st_4
      & (else_7_if_1_div_9cyc_st_4[0]) & (else_7_if_1_div_9cyc_st_4[1]) & (else_7_if_1_div_9cyc_st_4[2])
      & (~ (else_7_if_1_div_9cyc_st_4[3])));
  assign or_tmp_2166 = ~(main_stage_0_6 & (~ if_7_equal_svs_st_5) & else_7_equal_svs_st_5
      & (else_7_if_1_div_9cyc_st_5[0]) & (else_7_if_1_div_9cyc_st_5[1]) & (else_7_if_1_div_9cyc_st_5[2])
      & (~ (else_7_if_1_div_9cyc_st_5[3])));
  assign or_tmp_2173 = ~(main_stage_0_7 & (~ if_7_equal_svs_st_6) & else_7_equal_svs_st_6
      & (else_7_if_1_div_9cyc_st_6[0]) & (else_7_if_1_div_9cyc_st_6[1]) & (else_7_if_1_div_9cyc_st_6[2])
      & (~ (else_7_if_1_div_9cyc_st_6[3])));
  assign and_tmp_722 = or_tmp_2153 & or_tmp_2151;
  assign or_dcpl_935 = (~ (else_7_if_1_acc_tmp[3])) | (else_7_if_1_acc_tmp[0]) |
      (else_7_if_1_acc_tmp[2]);
  assign or_tmp_2231 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_9cyc_st_2[0]) | (else_7_if_1_div_9cyc_st_2[1]) | (else_7_if_1_div_9cyc_st_2[2]);
  assign or_tmp_2232 = (else_7_if_1_div_9cyc[0]) | (else_7_if_1_div_9cyc[1]) | (else_7_if_1_div_9cyc[2])
      | (~ (else_7_if_1_div_9cyc[3])) | (~ main_stage_0_2) | if_7_equal_svs_st_1;
  assign or_tmp_2233 = (~ (else_7_if_1_acc_tmp[3])) | (else_7_if_1_acc_tmp[2]) |
      (else_7_if_1_acc_tmp[1]) | (else_7_if_1_acc_tmp[0]) | (~ else_7_equal_tmp)
      | if_7_equal_tmp;
  assign mux_tmp_376 = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ or_tmp_2233)))
      , or_tmp_2233}, or_tmp_2232);
  assign or_tmp_2236 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | (~ else_7_equal_svs_st_3)
      | (else_7_if_1_div_9cyc_st_3[0]) | (else_7_if_1_div_9cyc_st_3[1]) | (else_7_if_1_div_9cyc_st_3[2]);
  assign or_tmp_2243 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | (~ else_7_equal_svs_st_4)
      | (else_7_if_1_div_9cyc_st_4[0]) | (else_7_if_1_div_9cyc_st_4[1]) | (else_7_if_1_div_9cyc_st_4[2]);
  assign mux_466_cse = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_3[3]) | (~ mux_460_cse)))
      , mux_460_cse}, or_tmp_2236);
  assign or_tmp_2252 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | (~ else_7_equal_svs_st_5)
      | (else_7_if_1_div_9cyc_st_5[0]) | (else_7_if_1_div_9cyc_st_5[1]) | (else_7_if_1_div_9cyc_st_5[2]);
  assign mux_471_cse = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_4[3]) | (~ mux_466_cse)))
      , mux_466_cse}, or_tmp_2243);
  assign and_tmp_755 = or_tmp_2233 & (or_tmp_2231 | (~ (else_7_if_1_div_9cyc_st_2[3])));
  assign mux_tmp_390 = MUX_s_1_2_2({(~(else_7_equal_svs_st_1 | (~ and_tmp_755)))
      , and_tmp_755}, or_tmp_2232);
  assign mux_tmp_391 = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_3[3]) | (~ mux_tmp_390)))
      , mux_tmp_390}, or_tmp_2236);
  assign mux_tmp_392 = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_4[3]) | (~ mux_tmp_391)))
      , mux_tmp_391}, or_tmp_2243);
  assign mux_476_cse = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_5[3]) | (~ mux_tmp_392)))
      , mux_tmp_392}, or_tmp_2252);
  assign mux_482_cse = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_6[3]) | (~ mux_476_cse)))
      , mux_476_cse}, (~ main_stage_0_7) | if_7_equal_svs_st_6 | (~ else_7_equal_svs_st_6)
      | (else_7_if_1_div_9cyc_st_6[0]) | (else_7_if_1_div_9cyc_st_6[1]) | (else_7_if_1_div_9cyc_st_6[2]));
  assign and_dcpl_4962 = ~((else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[0]));
  assign and_dcpl_4963 = and_dcpl_4962 & (~ (else_7_else_1_if_acc_tmp[2]));
  assign and_dcpl_4965 = ~(if_7_equal_tmp | else_7_equal_tmp);
  assign and_dcpl_4966 = and_dcpl_4965 & else_7_else_1_equal_tmp & (~ (else_7_else_1_if_acc_tmp[1]));
  assign and_dcpl_4968 = ~((else_7_else_1_if_div_9cyc[1]) | (else_7_else_1_if_div_9cyc[2]));
  assign and_dcpl_4969 = and_dcpl_4968 & (~ (else_7_else_1_if_div_9cyc[0]));
  assign and_dcpl_4971 = main_stage_0_2 & (~ else_7_equal_svs_st_1);
  assign and_dcpl_4972 = and_dcpl_4971 & else_7_else_1_equal_svs_1 & (~ (else_7_else_1_if_div_9cyc[3]));
  assign or_dcpl_944 = (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[0]);
  assign or_dcpl_945 = or_dcpl_944 | (else_7_else_1_if_acc_tmp[2]);
  assign or_dcpl_947 = if_7_equal_tmp | else_7_equal_tmp;
  assign or_dcpl_948 = or_dcpl_947 | (~ else_7_else_1_equal_tmp) | (else_7_else_1_if_acc_tmp[1]);
  assign and_dcpl_4981 = and_1994_cse & (~ else_7_equal_svs_st_2) & else_7_else_1_equal_svs_st_2;
  assign and_dcpl_4989 = and_1622_cse & (~ else_7_equal_svs_st_3) & else_7_else_1_equal_svs_st_3;
  assign or_tmp_2353 = (else_7_else_1_if_div_9cyc[0]) | (else_7_else_1_if_div_9cyc[1])
      | (else_7_else_1_if_div_9cyc[2]) | (else_7_else_1_if_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2354 = (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[2])
      | (else_7_else_1_if_acc_tmp[1]) | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2355 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_9cyc_st_2[0]) |
      (else_7_else_1_if_div_9cyc_st_2[1]) | (else_7_else_1_if_div_9cyc_st_2[2]) |
      (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_760 = or_tmp_2354 & or_tmp_2355;
  assign and_dcpl_4997 = and_1250_cse & (~ else_7_equal_svs_st_4) & else_7_else_1_equal_svs_st_4;
  assign or_tmp_2360 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_9cyc_st_3[0]) |
      (else_7_else_1_if_div_9cyc_st_3[1]) | (else_7_else_1_if_div_9cyc_st_3[2]) |
      (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_762 = or_tmp_2355 & or_tmp_2354 & or_tmp_2360;
  assign and_dcpl_5005 = and_878_cse & (~ else_7_equal_svs_st_5) & else_7_else_1_equal_svs_st_5;
  assign or_tmp_2363 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (else_7_else_1_if_div_9cyc_st_4[0]) |
      (else_7_else_1_if_div_9cyc_st_4[1]) | (else_7_else_1_if_div_9cyc_st_4[2]) |
      (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_763 = or_tmp_2355 & or_tmp_2354;
  assign and_tmp_765 = or_tmp_2363 & or_tmp_2360 & and_tmp_763;
  assign and_dcpl_5013 = and_506_cse & (~ else_7_equal_svs_st_6) & else_7_else_1_equal_svs_st_6;
  assign or_tmp_2369 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (else_7_else_1_if_div_9cyc_st_5[0]) |
      (else_7_else_1_if_div_9cyc_st_5[1]) | (else_7_else_1_if_div_9cyc_st_5[2]) |
      (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_769 = or_tmp_2369 & or_tmp_2363 & or_tmp_2360 & and_tmp_763;
  assign and_dcpl_5021 = and_dcpl_17 & (~ else_7_equal_svs_st_7) & else_7_else_1_equal_svs_st_7;
  assign or_tmp_2376 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (else_7_else_1_if_div_9cyc_st_6[0]) |
      (else_7_else_1_if_div_9cyc_st_6[1]) | (else_7_else_1_if_div_9cyc_st_6[2]) |
      (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_774 = or_tmp_2376 & or_tmp_2369 & or_tmp_2363 & or_tmp_2360 & and_tmp_763;
  assign and_tmp_780 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (else_7_else_1_if_div_9cyc_st_7[0]) |
      (else_7_else_1_if_div_9cyc_st_7[1]) | (else_7_else_1_if_div_9cyc_st_7[2]) |
      (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2354 & or_tmp_2376 & or_tmp_2369
      & or_tmp_2363 & or_tmp_2360 & or_tmp_2355;
  assign and_dcpl_5086 = (~ (else_7_else_1_if_acc_tmp[3])) & (else_7_else_1_if_acc_tmp[0]);
  assign and_dcpl_5087 = and_dcpl_5086 & (~ (else_7_else_1_if_acc_tmp[2]));
  assign or_dcpl_956 = (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[0]));
  assign or_dcpl_957 = or_dcpl_956 | (else_7_else_1_if_acc_tmp[2]);
  assign or_tmp_2433 = (~ (else_7_else_1_if_div_9cyc[0])) | (else_7_else_1_if_div_9cyc[1])
      | (else_7_else_1_if_div_9cyc[2]) | (else_7_else_1_if_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2434 = (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[2])
      | (else_7_else_1_if_acc_tmp[1]) | (~ (else_7_else_1_if_acc_tmp[0])) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2435 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (~ (else_7_else_1_if_div_9cyc_st_2[0]))
      | (else_7_else_1_if_div_9cyc_st_2[1]) | (else_7_else_1_if_div_9cyc_st_2[2])
      | (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_803 = or_tmp_2434 & or_tmp_2435;
  assign or_tmp_2440 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (~ (else_7_else_1_if_div_9cyc_st_3[0]))
      | (else_7_else_1_if_div_9cyc_st_3[1]) | (else_7_else_1_if_div_9cyc_st_3[2])
      | (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_805 = or_tmp_2435 & or_tmp_2434 & or_tmp_2440;
  assign or_tmp_2443 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (~ (else_7_else_1_if_div_9cyc_st_4[0]))
      | (else_7_else_1_if_div_9cyc_st_4[1]) | (else_7_else_1_if_div_9cyc_st_4[2])
      | (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_806 = or_tmp_2435 & or_tmp_2434;
  assign and_tmp_808 = or_tmp_2443 & or_tmp_2440 & and_tmp_806;
  assign or_tmp_2449 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (~ (else_7_else_1_if_div_9cyc_st_5[0]))
      | (else_7_else_1_if_div_9cyc_st_5[1]) | (else_7_else_1_if_div_9cyc_st_5[2])
      | (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_812 = or_tmp_2449 & or_tmp_2443 & or_tmp_2440 & and_tmp_806;
  assign or_tmp_2456 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (~ (else_7_else_1_if_div_9cyc_st_6[0]))
      | (else_7_else_1_if_div_9cyc_st_6[1]) | (else_7_else_1_if_div_9cyc_st_6[2])
      | (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_817 = or_tmp_2456 & or_tmp_2449 & or_tmp_2443 & or_tmp_2440 & and_tmp_806;
  assign and_tmp_823 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (~ (else_7_else_1_if_div_9cyc_st_7[0]))
      | (else_7_else_1_if_div_9cyc_st_7[1]) | (else_7_else_1_if_div_9cyc_st_7[2])
      | (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2434 & or_tmp_2456 & or_tmp_2449
      & or_tmp_2443 & or_tmp_2440 & or_tmp_2435;
  assign and_dcpl_5214 = and_dcpl_4965 & else_7_else_1_equal_tmp & (else_7_else_1_if_acc_tmp[1]);
  assign and_dcpl_5216 = (else_7_else_1_if_div_9cyc[1]) & (~ (else_7_else_1_if_div_9cyc[2]));
  assign or_dcpl_972 = or_dcpl_947 | (~(else_7_else_1_equal_tmp & (else_7_else_1_if_acc_tmp[1])));
  assign or_tmp_2513 = (else_7_else_1_if_div_9cyc[0]) | (~ (else_7_else_1_if_div_9cyc[1]))
      | (else_7_else_1_if_div_9cyc[2]) | (else_7_else_1_if_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2514 = (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[2])
      | (~ (else_7_else_1_if_acc_tmp[1])) | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2515 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_9cyc_st_2[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_2[1])) | (else_7_else_1_if_div_9cyc_st_2[2])
      | (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_846 = or_tmp_2514 & or_tmp_2515;
  assign or_tmp_2520 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_9cyc_st_3[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_3[1])) | (else_7_else_1_if_div_9cyc_st_3[2])
      | (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_848 = or_tmp_2515 & or_tmp_2514 & or_tmp_2520;
  assign or_tmp_2523 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (else_7_else_1_if_div_9cyc_st_4[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_4[1])) | (else_7_else_1_if_div_9cyc_st_4[2])
      | (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_849 = or_tmp_2515 & or_tmp_2514;
  assign and_tmp_851 = or_tmp_2523 & or_tmp_2520 & and_tmp_849;
  assign or_tmp_2529 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (else_7_else_1_if_div_9cyc_st_5[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_5[1])) | (else_7_else_1_if_div_9cyc_st_5[2])
      | (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_855 = or_tmp_2529 & or_tmp_2523 & or_tmp_2520 & and_tmp_849;
  assign or_tmp_2536 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (else_7_else_1_if_div_9cyc_st_6[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_6[1])) | (else_7_else_1_if_div_9cyc_st_6[2])
      | (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_860 = or_tmp_2536 & or_tmp_2529 & or_tmp_2523 & or_tmp_2520 & and_tmp_849;
  assign and_tmp_866 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (else_7_else_1_if_div_9cyc_st_7[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_7[1])) | (else_7_else_1_if_div_9cyc_st_7[2])
      | (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2514 & or_tmp_2536 & or_tmp_2529
      & or_tmp_2523 & or_tmp_2520 & or_tmp_2515;
  assign or_tmp_2593 = (~ (else_7_else_1_if_div_9cyc[0])) | (~ (else_7_else_1_if_div_9cyc[1]))
      | (else_7_else_1_if_div_9cyc[2]) | (else_7_else_1_if_div_9cyc[3]) | (~ main_stage_0_2)
      | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2594 = (else_7_else_1_if_acc_tmp[3]) | (else_7_else_1_if_acc_tmp[2])
      | (~ (else_7_else_1_if_acc_tmp[1])) | (~ (else_7_else_1_if_acc_tmp[0])) | (~
      else_7_else_1_equal_tmp) | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2595 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (~ (else_7_else_1_if_div_9cyc_st_2[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_2[1])) | (else_7_else_1_if_div_9cyc_st_2[2])
      | (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_889 = or_tmp_2594 & or_tmp_2595;
  assign or_tmp_2600 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (~ (else_7_else_1_if_div_9cyc_st_3[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_3[1])) | (else_7_else_1_if_div_9cyc_st_3[2])
      | (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_891 = or_tmp_2595 & or_tmp_2594 & or_tmp_2600;
  assign or_tmp_2603 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (~ (else_7_else_1_if_div_9cyc_st_4[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_4[1])) | (else_7_else_1_if_div_9cyc_st_4[2])
      | (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_892 = or_tmp_2595 & or_tmp_2594;
  assign and_tmp_894 = or_tmp_2603 & or_tmp_2600 & and_tmp_892;
  assign or_tmp_2609 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (~ (else_7_else_1_if_div_9cyc_st_5[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_5[1])) | (else_7_else_1_if_div_9cyc_st_5[2])
      | (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_898 = or_tmp_2609 & or_tmp_2603 & or_tmp_2600 & and_tmp_892;
  assign or_tmp_2616 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (~ (else_7_else_1_if_div_9cyc_st_6[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_6[1])) | (else_7_else_1_if_div_9cyc_st_6[2])
      | (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_903 = or_tmp_2616 & or_tmp_2609 & or_tmp_2603 & or_tmp_2600 & and_tmp_892;
  assign and_tmp_909 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (~ (else_7_else_1_if_div_9cyc_st_7[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_7[1])) | (else_7_else_1_if_div_9cyc_st_7[2])
      | (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2594 & or_tmp_2616 & or_tmp_2609
      & or_tmp_2603 & or_tmp_2600 & or_tmp_2595;
  assign and_dcpl_5459 = and_dcpl_4962 & (else_7_else_1_if_acc_tmp[2]);
  assign and_dcpl_5464 = (~ (else_7_else_1_if_div_9cyc[1])) & (else_7_else_1_if_div_9cyc[2]);
  assign or_dcpl_993 = or_dcpl_944 | (~ (else_7_else_1_if_acc_tmp[2]));
  assign or_tmp_2673 = (else_7_else_1_if_div_9cyc[0]) | (else_7_else_1_if_div_9cyc[1])
      | (~ (else_7_else_1_if_div_9cyc[2])) | (else_7_else_1_if_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2674 = (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[2]))
      | (else_7_else_1_if_acc_tmp[1]) | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2675 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_9cyc_st_2[0]) |
      (else_7_else_1_if_div_9cyc_st_2[1]) | (~ (else_7_else_1_if_div_9cyc_st_2[2]))
      | (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_932 = or_tmp_2674 & or_tmp_2675;
  assign or_tmp_2680 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_9cyc_st_3[0]) |
      (else_7_else_1_if_div_9cyc_st_3[1]) | (~ (else_7_else_1_if_div_9cyc_st_3[2]))
      | (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_934 = or_tmp_2675 & or_tmp_2674 & or_tmp_2680;
  assign or_tmp_2683 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (else_7_else_1_if_div_9cyc_st_4[0]) |
      (else_7_else_1_if_div_9cyc_st_4[1]) | (~ (else_7_else_1_if_div_9cyc_st_4[2]))
      | (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_935 = or_tmp_2675 & or_tmp_2674;
  assign and_tmp_937 = or_tmp_2683 & or_tmp_2680 & and_tmp_935;
  assign or_tmp_2689 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (else_7_else_1_if_div_9cyc_st_5[0]) |
      (else_7_else_1_if_div_9cyc_st_5[1]) | (~ (else_7_else_1_if_div_9cyc_st_5[2]))
      | (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_941 = or_tmp_2689 & or_tmp_2683 & or_tmp_2680 & and_tmp_935;
  assign or_tmp_2696 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (else_7_else_1_if_div_9cyc_st_6[0]) |
      (else_7_else_1_if_div_9cyc_st_6[1]) | (~ (else_7_else_1_if_div_9cyc_st_6[2]))
      | (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_946 = or_tmp_2696 & or_tmp_2689 & or_tmp_2683 & or_tmp_2680 & and_tmp_935;
  assign and_tmp_952 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (else_7_else_1_if_div_9cyc_st_7[0]) |
      (else_7_else_1_if_div_9cyc_st_7[1]) | (~ (else_7_else_1_if_div_9cyc_st_7[2]))
      | (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2674 & or_tmp_2696 & or_tmp_2689
      & or_tmp_2683 & or_tmp_2680 & or_tmp_2675;
  assign and_dcpl_5583 = and_dcpl_5086 & (else_7_else_1_if_acc_tmp[2]);
  assign or_dcpl_1005 = or_dcpl_956 | (~ (else_7_else_1_if_acc_tmp[2]));
  assign or_tmp_2753 = (~ (else_7_else_1_if_div_9cyc[0])) | (else_7_else_1_if_div_9cyc[1])
      | (~ (else_7_else_1_if_div_9cyc[2])) | (else_7_else_1_if_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2754 = (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[2]))
      | (else_7_else_1_if_acc_tmp[1]) | (~ (else_7_else_1_if_acc_tmp[0])) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2755 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (~ (else_7_else_1_if_div_9cyc_st_2[0]))
      | (else_7_else_1_if_div_9cyc_st_2[1]) | (~ (else_7_else_1_if_div_9cyc_st_2[2]))
      | (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_975 = or_tmp_2754 & or_tmp_2755;
  assign or_tmp_2760 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (~ (else_7_else_1_if_div_9cyc_st_3[0]))
      | (else_7_else_1_if_div_9cyc_st_3[1]) | (~ (else_7_else_1_if_div_9cyc_st_3[2]))
      | (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_977 = or_tmp_2755 & or_tmp_2754 & or_tmp_2760;
  assign or_tmp_2763 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (~ (else_7_else_1_if_div_9cyc_st_4[0]))
      | (else_7_else_1_if_div_9cyc_st_4[1]) | (~ (else_7_else_1_if_div_9cyc_st_4[2]))
      | (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_978 = or_tmp_2755 & or_tmp_2754;
  assign and_tmp_980 = or_tmp_2763 & or_tmp_2760 & and_tmp_978;
  assign or_tmp_2769 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (~ (else_7_else_1_if_div_9cyc_st_5[0]))
      | (else_7_else_1_if_div_9cyc_st_5[1]) | (~ (else_7_else_1_if_div_9cyc_st_5[2]))
      | (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_984 = or_tmp_2769 & or_tmp_2763 & or_tmp_2760 & and_tmp_978;
  assign or_tmp_2776 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (~ (else_7_else_1_if_div_9cyc_st_6[0]))
      | (else_7_else_1_if_div_9cyc_st_6[1]) | (~ (else_7_else_1_if_div_9cyc_st_6[2]))
      | (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_989 = or_tmp_2776 & or_tmp_2769 & or_tmp_2763 & or_tmp_2760 & and_tmp_978;
  assign and_tmp_995 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (~ (else_7_else_1_if_div_9cyc_st_7[0]))
      | (else_7_else_1_if_div_9cyc_st_7[1]) | (~ (else_7_else_1_if_div_9cyc_st_7[2]))
      | (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2754 & or_tmp_2776 & or_tmp_2769
      & or_tmp_2763 & or_tmp_2760 & or_tmp_2755;
  assign and_dcpl_5712 = (else_7_else_1_if_div_9cyc[1]) & (else_7_else_1_if_div_9cyc[2]);
  assign or_tmp_2833 = (else_7_else_1_if_div_9cyc[0]) | (~ (else_7_else_1_if_div_9cyc[1]))
      | (~ (else_7_else_1_if_div_9cyc[2])) | (else_7_else_1_if_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2834 = (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[2]))
      | (~ (else_7_else_1_if_acc_tmp[1])) | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2835 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_9cyc_st_2[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_2[1])) | (~ (else_7_else_1_if_div_9cyc_st_2[2]))
      | (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_1018 = or_tmp_2834 & or_tmp_2835;
  assign or_tmp_2840 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_9cyc_st_3[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_3[1])) | (~ (else_7_else_1_if_div_9cyc_st_3[2]))
      | (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_1020 = or_tmp_2835 & or_tmp_2834 & or_tmp_2840;
  assign or_tmp_2843 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (else_7_else_1_if_div_9cyc_st_4[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_4[1])) | (~ (else_7_else_1_if_div_9cyc_st_4[2]))
      | (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_1021 = or_tmp_2835 & or_tmp_2834;
  assign and_tmp_1023 = or_tmp_2843 & or_tmp_2840 & and_tmp_1021;
  assign or_tmp_2849 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (else_7_else_1_if_div_9cyc_st_5[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_5[1])) | (~ (else_7_else_1_if_div_9cyc_st_5[2]))
      | (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_1027 = or_tmp_2849 & or_tmp_2843 & or_tmp_2840 & and_tmp_1021;
  assign or_tmp_2856 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (else_7_else_1_if_div_9cyc_st_6[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_6[1])) | (~ (else_7_else_1_if_div_9cyc_st_6[2]))
      | (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_1032 = or_tmp_2856 & or_tmp_2849 & or_tmp_2843 & or_tmp_2840 & and_tmp_1021;
  assign and_tmp_1038 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (else_7_else_1_if_div_9cyc_st_7[0]) |
      (~ (else_7_else_1_if_div_9cyc_st_7[1])) | (~ (else_7_else_1_if_div_9cyc_st_7[2]))
      | (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2834 & or_tmp_2856 & or_tmp_2849
      & or_tmp_2843 & or_tmp_2840 & or_tmp_2835;
  assign or_tmp_2913 = (~ (else_7_else_1_if_div_9cyc[0])) | (~ (else_7_else_1_if_div_9cyc[1]))
      | (~ (else_7_else_1_if_div_9cyc[2])) | (else_7_else_1_if_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2914 = (else_7_else_1_if_acc_tmp[3]) | (~ (else_7_else_1_if_acc_tmp[2]))
      | (~ (else_7_else_1_if_acc_tmp[1])) | (~ (else_7_else_1_if_acc_tmp[0])) | (~
      else_7_else_1_equal_tmp) | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2915 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (~ (else_7_else_1_if_div_9cyc_st_2[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_2[1])) | (~ (else_7_else_1_if_div_9cyc_st_2[2]))
      | (else_7_else_1_if_div_9cyc_st_2[3]);
  assign and_tmp_1061 = or_tmp_2914 & or_tmp_2915;
  assign or_tmp_2920 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (~ (else_7_else_1_if_div_9cyc_st_3[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_3[1])) | (~ (else_7_else_1_if_div_9cyc_st_3[2]))
      | (else_7_else_1_if_div_9cyc_st_3[3]);
  assign and_tmp_1063 = or_tmp_2915 & or_tmp_2914 & or_tmp_2920;
  assign or_tmp_2923 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (~ (else_7_else_1_if_div_9cyc_st_4[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_4[1])) | (~ (else_7_else_1_if_div_9cyc_st_4[2]))
      | (else_7_else_1_if_div_9cyc_st_4[3]);
  assign and_tmp_1064 = or_tmp_2915 & or_tmp_2914;
  assign and_tmp_1066 = or_tmp_2923 & or_tmp_2920 & and_tmp_1064;
  assign or_tmp_2929 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (~ (else_7_else_1_if_div_9cyc_st_5[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_5[1])) | (~ (else_7_else_1_if_div_9cyc_st_5[2]))
      | (else_7_else_1_if_div_9cyc_st_5[3]);
  assign and_tmp_1070 = or_tmp_2929 & or_tmp_2923 & or_tmp_2920 & and_tmp_1064;
  assign or_tmp_2936 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (~ (else_7_else_1_if_div_9cyc_st_6[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_6[1])) | (~ (else_7_else_1_if_div_9cyc_st_6[2]))
      | (else_7_else_1_if_div_9cyc_st_6[3]);
  assign and_tmp_1075 = or_tmp_2936 & or_tmp_2929 & or_tmp_2923 & or_tmp_2920 & and_tmp_1064;
  assign and_tmp_1081 = ((~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (~ (else_7_else_1_if_div_9cyc_st_7[0]))
      | (~ (else_7_else_1_if_div_9cyc_st_7[1])) | (~ (else_7_else_1_if_div_9cyc_st_7[2]))
      | (else_7_else_1_if_div_9cyc_st_7[3])) & or_tmp_2914 & or_tmp_2936 & or_tmp_2929
      & or_tmp_2923 & or_tmp_2920 & or_tmp_2915;
  assign or_dcpl_1041 = (~ (else_7_else_1_if_acc_tmp[3])) | (else_7_else_1_if_acc_tmp[0])
      | (else_7_else_1_if_acc_tmp[2]);
  assign or_tmp_2993 = (else_7_else_1_if_div_9cyc[0]) | (else_7_else_1_if_div_9cyc[1])
      | (else_7_else_1_if_div_9cyc[2]) | (~ (else_7_else_1_if_div_9cyc[3])) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1;
  assign or_tmp_2994 = (~ (else_7_else_1_if_acc_tmp[3])) | (else_7_else_1_if_acc_tmp[2])
      | (else_7_else_1_if_acc_tmp[1]) | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp)
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_2995 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_9cyc_st_2[0]) |
      (else_7_else_1_if_div_9cyc_st_2[1]) | (else_7_else_1_if_div_9cyc_st_2[2]);
  assign or_tmp_2996 = or_tmp_2995 | (~ (else_7_else_1_if_div_9cyc_st_2[3]));
  assign and_tmp_1104 = or_tmp_2994 & or_tmp_2996;
  assign or_tmp_3001 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_9cyc_st_3[0]) |
      (else_7_else_1_if_div_9cyc_st_3[1]) | (else_7_else_1_if_div_9cyc_st_3[2]);
  assign and_tmp_1105 = or_tmp_2994 & (or_tmp_3001 | (~ (else_7_else_1_if_div_9cyc_st_3[3])));
  assign mux_tmp_523 = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_2[3]) | (~ and_tmp_1105)))
      , and_tmp_1105}, or_tmp_2995);
  assign or_tmp_3006 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | (~ else_7_else_1_equal_svs_st_4) | (else_7_else_1_if_div_9cyc_st_4[0]) |
      (else_7_else_1_if_div_9cyc_st_4[1]) | (else_7_else_1_if_div_9cyc_st_4[2]);
  assign mux_tmp_525 = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_2[3]) | (~ or_tmp_2994)))
      , or_tmp_2994}, or_tmp_2995);
  assign mux_tmp_526 = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_3[3]) | (~ mux_tmp_525)))
      , mux_tmp_525}, or_tmp_3001);
  assign mux_610_cse = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_4[3]) | (~ mux_tmp_526)))
      , mux_tmp_526}, or_tmp_3006);
  assign or_tmp_3015 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | (~ else_7_else_1_equal_svs_st_5) | (else_7_else_1_if_div_9cyc_st_5[0]) |
      (else_7_else_1_if_div_9cyc_st_5[1]) | (else_7_else_1_if_div_9cyc_st_5[2]);
  assign mux_615_cse = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_5[3]) | (~ mux_610_cse)))
      , mux_610_cse}, or_tmp_3015);
  assign or_tmp_3026 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | (~ else_7_else_1_equal_svs_st_6) | (else_7_else_1_if_div_9cyc_st_6[0]) |
      (else_7_else_1_if_div_9cyc_st_6[1]) | (else_7_else_1_if_div_9cyc_st_6[2]);
  assign mux_621_cse = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_6[3]) | (~ mux_615_cse)))
      , mux_615_cse}, or_tmp_3026);
  assign mux_tmp_540 = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_3[3]) | (~ or_tmp_2996)))
      , or_tmp_2996}, or_tmp_3001);
  assign mux_tmp_541 = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_4[3]) | (~ mux_tmp_540)))
      , mux_tmp_540}, or_tmp_3006);
  assign mux_tmp_542 = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_5[3]) | (~ mux_tmp_541)))
      , mux_tmp_541}, or_tmp_3015);
  assign mux_626_nl = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_6[3]) | (~ mux_tmp_542)))
      , mux_tmp_542}, or_tmp_3026);
  assign and_tmp_1106 = or_tmp_2994 & (mux_626_nl);
  assign mux_627_cse = MUX_s_1_2_2({(~((else_7_else_1_if_div_9cyc_st_7[3]) | (~ and_tmp_1106)))
      , and_tmp_1106}, (~ main_stage_0_8) | if_7_equal_svs_st_7 | else_7_equal_svs_st_7
      | (~ else_7_else_1_equal_svs_st_7) | (else_7_else_1_if_div_9cyc_st_7[0]) |
      (else_7_else_1_if_div_9cyc_st_7[1]) | (else_7_else_1_if_div_9cyc_st_7[2]));
  assign and_dcpl_6078 = ~((else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[0]));
  assign and_dcpl_6079 = and_dcpl_6078 & (~ (else_7_else_1_else_acc_tmp[2]));
  assign and_dcpl_6082 = and_dcpl_4965 & (~(else_7_else_1_equal_tmp | (else_7_else_1_else_acc_tmp[1])));
  assign and_dcpl_6084 = ~((else_7_else_1_else_div_9cyc[3]) | (else_7_else_1_else_div_9cyc[1]));
  assign and_dcpl_6085 = and_dcpl_6084 & (~ (else_7_else_1_else_div_9cyc[0]));
  assign and_dcpl_6088 = and_dcpl_4971 & (~(else_7_else_1_equal_svs_1 | (else_7_else_1_else_div_9cyc[2])));
  assign or_dcpl_1052 = (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[0]);
  assign or_dcpl_1053 = or_dcpl_1052 | (else_7_else_1_else_acc_tmp[2]);
  assign or_dcpl_1056 = or_dcpl_947 | else_7_else_1_equal_tmp | (else_7_else_1_else_acc_tmp[1]);
  assign or_tmp_3115 = (else_7_else_1_else_div_9cyc[0]) | (else_7_else_1_else_div_9cyc[1])
      | (else_7_else_1_else_div_9cyc[2]) | (else_7_else_1_else_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3116 = (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[2])
      | (else_7_else_1_else_acc_tmp[1]) | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3117 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_9cyc_st_2[0]) | (else_7_else_1_else_div_9cyc_st_2[1])
      | (else_7_else_1_else_div_9cyc_st_2[2]) | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3121 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_9cyc_st_3[0]) | (else_7_else_1_else_div_9cyc_st_3[1])
      | (else_7_else_1_else_div_9cyc_st_3[2]) | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3123 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (else_7_else_1_else_div_9cyc_st_4[0]) | (else_7_else_1_else_div_9cyc_st_4[1])
      | (else_7_else_1_else_div_9cyc_st_4[2]) | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1116 = or_tmp_3117 & or_tmp_3116;
  assign or_tmp_3128 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (else_7_else_1_else_div_9cyc_st_5[0]) | (else_7_else_1_else_div_9cyc_st_5[1])
      | (else_7_else_1_else_div_9cyc_st_5[2]) | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3134 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (else_7_else_1_else_div_9cyc_st_6[0]) | (else_7_else_1_else_div_9cyc_st_6[1])
      | (else_7_else_1_else_div_9cyc_st_6[2]) | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign and_dcpl_6202 = (~ (else_7_else_1_else_acc_tmp[3])) & (else_7_else_1_else_acc_tmp[0]);
  assign and_dcpl_6203 = and_dcpl_6202 & (~ (else_7_else_1_else_acc_tmp[2]));
  assign and_dcpl_6209 = and_dcpl_6084 & (else_7_else_1_else_div_9cyc[0]);
  assign or_dcpl_1064 = (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[0]));
  assign or_dcpl_1065 = or_dcpl_1064 | (else_7_else_1_else_acc_tmp[2]);
  assign or_tmp_3183 = (~ (else_7_else_1_else_div_9cyc[0])) | (else_7_else_1_else_div_9cyc[1])
      | (else_7_else_1_else_div_9cyc[2]) | (else_7_else_1_else_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3184 = (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[2])
      | (else_7_else_1_else_acc_tmp[1]) | (~ (else_7_else_1_else_acc_tmp[0])) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3185 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (~ (else_7_else_1_else_div_9cyc_st_2[0]))
      | (else_7_else_1_else_div_9cyc_st_2[1]) | (else_7_else_1_else_div_9cyc_st_2[2])
      | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3189 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (~ (else_7_else_1_else_div_9cyc_st_3[0]))
      | (else_7_else_1_else_div_9cyc_st_3[1]) | (else_7_else_1_else_div_9cyc_st_3[2])
      | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3191 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (~ (else_7_else_1_else_div_9cyc_st_4[0]))
      | (else_7_else_1_else_div_9cyc_st_4[1]) | (else_7_else_1_else_div_9cyc_st_4[2])
      | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1171 = or_tmp_3185 & or_tmp_3184;
  assign or_tmp_3196 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (~ (else_7_else_1_else_div_9cyc_st_5[0]))
      | (else_7_else_1_else_div_9cyc_st_5[1]) | (else_7_else_1_else_div_9cyc_st_5[2])
      | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3202 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (~ (else_7_else_1_else_div_9cyc_st_6[0]))
      | (else_7_else_1_else_div_9cyc_st_6[1]) | (else_7_else_1_else_div_9cyc_st_6[2])
      | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign and_dcpl_6330 = and_dcpl_4965 & (~ else_7_else_1_equal_tmp) & (else_7_else_1_else_acc_tmp[1]);
  assign and_dcpl_6332 = (~ (else_7_else_1_else_div_9cyc[3])) & (else_7_else_1_else_div_9cyc[1]);
  assign and_dcpl_6333 = and_dcpl_6332 & (~ (else_7_else_1_else_div_9cyc[0]));
  assign or_dcpl_1080 = or_dcpl_947 | else_7_else_1_equal_tmp | (~ (else_7_else_1_else_acc_tmp[1]));
  assign or_tmp_3251 = (else_7_else_1_else_div_9cyc[0]) | (~ (else_7_else_1_else_div_9cyc[1]))
      | (else_7_else_1_else_div_9cyc[2]) | (else_7_else_1_else_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3252 = (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[2])
      | (~ (else_7_else_1_else_acc_tmp[1])) | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3253 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_9cyc_st_2[0]) | (~
      (else_7_else_1_else_div_9cyc_st_2[1])) | (else_7_else_1_else_div_9cyc_st_2[2])
      | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3257 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_9cyc_st_3[0]) | (~
      (else_7_else_1_else_div_9cyc_st_3[1])) | (else_7_else_1_else_div_9cyc_st_3[2])
      | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3259 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (else_7_else_1_else_div_9cyc_st_4[0]) | (~
      (else_7_else_1_else_div_9cyc_st_4[1])) | (else_7_else_1_else_div_9cyc_st_4[2])
      | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1226 = or_tmp_3253 & or_tmp_3252;
  assign or_tmp_3264 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (else_7_else_1_else_div_9cyc_st_5[0]) | (~
      (else_7_else_1_else_div_9cyc_st_5[1])) | (else_7_else_1_else_div_9cyc_st_5[2])
      | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3270 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (else_7_else_1_else_div_9cyc_st_6[0]) | (~
      (else_7_else_1_else_div_9cyc_st_6[1])) | (else_7_else_1_else_div_9cyc_st_6[2])
      | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign and_dcpl_6457 = and_dcpl_6332 & (else_7_else_1_else_div_9cyc[0]);
  assign or_tmp_3319 = (~ (else_7_else_1_else_div_9cyc[0])) | (~ (else_7_else_1_else_div_9cyc[1]))
      | (else_7_else_1_else_div_9cyc[2]) | (else_7_else_1_else_div_9cyc[3]) | (~
      main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3320 = (else_7_else_1_else_acc_tmp[3]) | (else_7_else_1_else_acc_tmp[2])
      | (~ (else_7_else_1_else_acc_tmp[1])) | (~ (else_7_else_1_else_acc_tmp[0]))
      | else_7_else_1_equal_tmp | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3321 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (~ (else_7_else_1_else_div_9cyc_st_2[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_2[1])) | (else_7_else_1_else_div_9cyc_st_2[2])
      | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3325 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (~ (else_7_else_1_else_div_9cyc_st_3[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_3[1])) | (else_7_else_1_else_div_9cyc_st_3[2])
      | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3327 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (~ (else_7_else_1_else_div_9cyc_st_4[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_4[1])) | (else_7_else_1_else_div_9cyc_st_4[2])
      | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1281 = or_tmp_3321 & or_tmp_3320;
  assign or_tmp_3332 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (~ (else_7_else_1_else_div_9cyc_st_5[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_5[1])) | (else_7_else_1_else_div_9cyc_st_5[2])
      | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3338 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (~ (else_7_else_1_else_div_9cyc_st_6[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_6[1])) | (else_7_else_1_else_div_9cyc_st_6[2])
      | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign and_dcpl_6575 = and_dcpl_6078 & (else_7_else_1_else_acc_tmp[2]);
  assign and_dcpl_6584 = and_dcpl_4971 & (~ else_7_else_1_equal_svs_1) & (else_7_else_1_else_div_9cyc[2]);
  assign or_dcpl_1101 = or_dcpl_1052 | (~ (else_7_else_1_else_acc_tmp[2]));
  assign or_tmp_3387 = (else_7_else_1_else_div_9cyc[0]) | (else_7_else_1_else_div_9cyc[1])
      | (~ (else_7_else_1_else_div_9cyc[2])) | (else_7_else_1_else_div_9cyc[3]) |
      (~ main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3388 = (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[2]))
      | (else_7_else_1_else_acc_tmp[1]) | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3389 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_9cyc_st_2[0]) | (else_7_else_1_else_div_9cyc_st_2[1])
      | (~ (else_7_else_1_else_div_9cyc_st_2[2])) | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3393 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_9cyc_st_3[0]) | (else_7_else_1_else_div_9cyc_st_3[1])
      | (~ (else_7_else_1_else_div_9cyc_st_3[2])) | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3395 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (else_7_else_1_else_div_9cyc_st_4[0]) | (else_7_else_1_else_div_9cyc_st_4[1])
      | (~ (else_7_else_1_else_div_9cyc_st_4[2])) | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1336 = or_tmp_3389 & or_tmp_3388;
  assign or_tmp_3400 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (else_7_else_1_else_div_9cyc_st_5[0]) | (else_7_else_1_else_div_9cyc_st_5[1])
      | (~ (else_7_else_1_else_div_9cyc_st_5[2])) | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3406 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (else_7_else_1_else_div_9cyc_st_6[0]) | (else_7_else_1_else_div_9cyc_st_6[1])
      | (~ (else_7_else_1_else_div_9cyc_st_6[2])) | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign and_dcpl_6699 = and_dcpl_6202 & (else_7_else_1_else_acc_tmp[2]);
  assign or_dcpl_1113 = or_dcpl_1064 | (~ (else_7_else_1_else_acc_tmp[2]));
  assign or_tmp_3455 = (~ (else_7_else_1_else_div_9cyc[0])) | (else_7_else_1_else_div_9cyc[1])
      | (~ (else_7_else_1_else_div_9cyc[2])) | (else_7_else_1_else_div_9cyc[3]) |
      (~ main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3456 = (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[2]))
      | (else_7_else_1_else_acc_tmp[1]) | (~ (else_7_else_1_else_acc_tmp[0])) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3457 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (~ (else_7_else_1_else_div_9cyc_st_2[0]))
      | (else_7_else_1_else_div_9cyc_st_2[1]) | (~ (else_7_else_1_else_div_9cyc_st_2[2]))
      | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3461 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (~ (else_7_else_1_else_div_9cyc_st_3[0]))
      | (else_7_else_1_else_div_9cyc_st_3[1]) | (~ (else_7_else_1_else_div_9cyc_st_3[2]))
      | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3463 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (~ (else_7_else_1_else_div_9cyc_st_4[0]))
      | (else_7_else_1_else_div_9cyc_st_4[1]) | (~ (else_7_else_1_else_div_9cyc_st_4[2]))
      | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1391 = or_tmp_3457 & or_tmp_3456;
  assign or_tmp_3468 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (~ (else_7_else_1_else_div_9cyc_st_5[0]))
      | (else_7_else_1_else_div_9cyc_st_5[1]) | (~ (else_7_else_1_else_div_9cyc_st_5[2]))
      | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3474 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (~ (else_7_else_1_else_div_9cyc_st_6[0]))
      | (else_7_else_1_else_div_9cyc_st_6[1]) | (~ (else_7_else_1_else_div_9cyc_st_6[2]))
      | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign or_tmp_3523 = (else_7_else_1_else_div_9cyc[0]) | (~ (else_7_else_1_else_div_9cyc[1]))
      | (~ (else_7_else_1_else_div_9cyc[2])) | (else_7_else_1_else_div_9cyc[3]) |
      (~ main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3524 = (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[2]))
      | (~ (else_7_else_1_else_acc_tmp[1])) | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3525 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_9cyc_st_2[0]) | (~
      (else_7_else_1_else_div_9cyc_st_2[1])) | (~ (else_7_else_1_else_div_9cyc_st_2[2]))
      | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3529 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_9cyc_st_3[0]) | (~
      (else_7_else_1_else_div_9cyc_st_3[1])) | (~ (else_7_else_1_else_div_9cyc_st_3[2]))
      | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3531 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (else_7_else_1_else_div_9cyc_st_4[0]) | (~
      (else_7_else_1_else_div_9cyc_st_4[1])) | (~ (else_7_else_1_else_div_9cyc_st_4[2]))
      | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1446 = or_tmp_3525 & or_tmp_3524;
  assign or_tmp_3536 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (else_7_else_1_else_div_9cyc_st_5[0]) | (~
      (else_7_else_1_else_div_9cyc_st_5[1])) | (~ (else_7_else_1_else_div_9cyc_st_5[2]))
      | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3542 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (else_7_else_1_else_div_9cyc_st_6[0]) | (~
      (else_7_else_1_else_div_9cyc_st_6[1])) | (~ (else_7_else_1_else_div_9cyc_st_6[2]))
      | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign or_tmp_3591 = (~ (else_7_else_1_else_div_9cyc[0])) | (~ (else_7_else_1_else_div_9cyc[1]))
      | (~ (else_7_else_1_else_div_9cyc[2])) | (else_7_else_1_else_div_9cyc[3]) |
      (~ main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3592 = (else_7_else_1_else_acc_tmp[3]) | (~ (else_7_else_1_else_acc_tmp[2]))
      | (~ (else_7_else_1_else_acc_tmp[1])) | (~ (else_7_else_1_else_acc_tmp[0]))
      | else_7_else_1_equal_tmp | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3593 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (~ (else_7_else_1_else_div_9cyc_st_2[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_2[1])) | (~ (else_7_else_1_else_div_9cyc_st_2[2]))
      | (else_7_else_1_else_div_9cyc_st_2[3]);
  assign or_tmp_3597 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (~ (else_7_else_1_else_div_9cyc_st_3[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_3[1])) | (~ (else_7_else_1_else_div_9cyc_st_3[2]))
      | (else_7_else_1_else_div_9cyc_st_3[3]);
  assign or_tmp_3599 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (~ (else_7_else_1_else_div_9cyc_st_4[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_4[1])) | (~ (else_7_else_1_else_div_9cyc_st_4[2]))
      | (else_7_else_1_else_div_9cyc_st_4[3]);
  assign and_tmp_1501 = or_tmp_3593 & or_tmp_3592;
  assign or_tmp_3604 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (~ (else_7_else_1_else_div_9cyc_st_5[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_5[1])) | (~ (else_7_else_1_else_div_9cyc_st_5[2]))
      | (else_7_else_1_else_div_9cyc_st_5[3]);
  assign or_tmp_3610 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (~ (else_7_else_1_else_div_9cyc_st_6[0]))
      | (~ (else_7_else_1_else_div_9cyc_st_6[1])) | (~ (else_7_else_1_else_div_9cyc_st_6[2]))
      | (else_7_else_1_else_div_9cyc_st_6[3]);
  assign or_dcpl_1149 = (~ (else_7_else_1_else_acc_tmp[3])) | (else_7_else_1_else_acc_tmp[0])
      | (else_7_else_1_else_acc_tmp[2]);
  assign or_tmp_3659 = (else_7_else_1_else_div_9cyc[0]) | (else_7_else_1_else_div_9cyc[1])
      | (else_7_else_1_else_div_9cyc[2]) | (~ (else_7_else_1_else_div_9cyc[3])) |
      (~ main_stage_0_2) | if_7_equal_svs_st_1 | else_7_equal_svs_st_1 | else_7_else_1_equal_svs_1;
  assign or_tmp_3660 = (~ (else_7_else_1_else_acc_tmp[3])) | (else_7_else_1_else_acc_tmp[2])
      | (else_7_else_1_else_acc_tmp[1]) | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp
      | else_7_equal_tmp | if_7_equal_tmp;
  assign or_tmp_3661 = (~ main_stage_0_3) | if_7_equal_svs_st_2 | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_9cyc_st_2[0]) | (else_7_else_1_else_div_9cyc_st_2[1])
      | (else_7_else_1_else_div_9cyc_st_2[2]);
  assign or_tmp_3662 = or_tmp_3661 | (~ (else_7_else_1_else_div_9cyc_st_2[3]));
  assign or_tmp_3666 = (~ main_stage_0_4) | if_7_equal_svs_st_3 | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_9cyc_st_3[0]) | (else_7_else_1_else_div_9cyc_st_3[1])
      | (else_7_else_1_else_div_9cyc_st_3[2]);
  assign and_tmp_1553 = or_tmp_3660 & (or_tmp_3666 | (~ (else_7_else_1_else_div_9cyc_st_3[3])));
  assign or_tmp_3670 = (~ main_stage_0_5) | if_7_equal_svs_st_4 | else_7_equal_svs_st_4
      | else_7_else_1_equal_svs_st_4 | (else_7_else_1_else_div_9cyc_st_4[0]) | (else_7_else_1_else_div_9cyc_st_4[1])
      | (else_7_else_1_else_div_9cyc_st_4[2]);
  assign mux_tmp_571 = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_2[3]) | (~
      or_tmp_3660))) , or_tmp_3660}, or_tmp_3661);
  assign mux_tmp_572 = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_3[3]) | (~
      mux_tmp_571))) , mux_tmp_571}, or_tmp_3666);
  assign or_tmp_3678 = (~ main_stage_0_6) | if_7_equal_svs_st_5 | else_7_equal_svs_st_5
      | else_7_else_1_equal_svs_st_5 | (else_7_else_1_else_div_9cyc_st_5[0]) | (else_7_else_1_else_div_9cyc_st_5[1])
      | (else_7_else_1_else_div_9cyc_st_5[2]);
  assign mux_659_cse = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_4[3]) | (~
      mux_tmp_572))) , mux_tmp_572}, or_tmp_3670);
  assign or_tmp_3688 = (~ main_stage_0_7) | if_7_equal_svs_st_6 | else_7_equal_svs_st_6
      | else_7_else_1_equal_svs_st_6 | (else_7_else_1_else_div_9cyc_st_6[0]) | (else_7_else_1_else_div_9cyc_st_6[1])
      | (else_7_else_1_else_div_9cyc_st_6[2]);
  assign mux_664_cse = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_5[3]) | (~
      mux_659_cse))) , mux_659_cse}, or_tmp_3678);
  assign mux_tmp_583 = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_3[3]) | (~
      or_tmp_3662))) , or_tmp_3662}, or_tmp_3666);
  assign mux_tmp_584 = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_4[3]) | (~
      mux_tmp_583))) , mux_tmp_583}, or_tmp_3670);
  assign mux_tmp_585 = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_5[3]) | (~
      mux_tmp_584))) , mux_tmp_584}, or_tmp_3678);
  assign mux_669_nl = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_6[3]) | (~
      mux_tmp_585))) , mux_tmp_585}, or_tmp_3688);
  assign and_8701_cse = or_tmp_3660 & (mux_669_nl);
  assign or_dcpl_1160 = (else_7_if_acc_tmp[1]) | (else_7_if_acc_tmp[0]);
  assign or_dcpl_1161 = if_7_equal_tmp | (else_7_if_acc_tmp[3]);
  assign or_dcpl_1162 = or_dcpl_1161 | (else_7_if_acc_tmp[2]);
  assign or_dcpl_1170 = (else_7_if_acc_tmp[1]) | (~ (else_7_if_acc_tmp[0]));
  assign or_dcpl_1180 = (~ (else_7_if_acc_tmp[1])) | (else_7_if_acc_tmp[0]);
  assign or_dcpl_1190 = ~((else_7_if_acc_tmp[1]) & (else_7_if_acc_tmp[0]));
  assign or_dcpl_1202 = or_dcpl_1161 | (~ (else_7_if_acc_tmp[2]));
  assign mux_93_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp))) , and_tmp}, or_tmp_9);
  assign and_3172_cse = (mux_93_nl) & and_dcpl_3158 & and_dcpl_3156;
  assign mux_94_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_1))) , and_tmp_1}, or_tmp_9);
  assign and_3180_cse = or_tmp_15 & (mux_94_nl) & and_dcpl_3164 & and_dcpl_3162;
  assign and_3189_cse = or_tmp_23 & or_626_cse & or_628_cse & mux_95_cse & and_dcpl_3170
      & and_dcpl_3168;
  assign and_3199_cse = or_tmp_33 & ((~ or_tmp_34) | (else_7_if_div_9cyc_st_4[3])
      | (else_7_if_div_9cyc_st_4[2]) | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_626_cse & or_628_cse & mux_95_cse
      & and_dcpl_3176 & and_dcpl_3174;
  assign mux_100_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_14))) , and_tmp_14},
      or_630_cse);
  assign and_3221_cse = ((~ or_tmp_60) | (else_7_if_div_9cyc_st_6[3]) | (else_7_if_div_9cyc_st_6[2])
      | (else_7_if_div_9cyc_st_6[1]) | (else_7_if_div_9cyc_st_6[0]) | (~ main_stage_0_7)
      | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (else_7_if_div_9cyc_st_5[3]) | (else_7_if_div_9cyc_st_5[2])
      | (else_7_if_div_9cyc_st_5[1]) | (else_7_if_div_9cyc_st_5[0]) | (~ main_stage_0_6)
      | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_626_cse & or_628_cse & (mux_100_nl) & and_dcpl_3188
      & and_dcpl_3186;
  assign mux_98_nl = MUX_s_1_2_2({and_3207_cse , (~(or_tmp_58 | (~ and_3207_cse)))},
      main_stage_0_6);
  assign mux_99_nl = MUX_s_1_2_2({(mux_98_nl) , and_3207_cse}, or_tmp_46);
  assign and_3209_cse = or_tmp_45 & (mux_99_nl) & and_dcpl_3182 & and_dcpl_3180;
  assign mux_106_cse = MUX_s_1_2_2({(~(or_tmp_94 | (~ mux_105_cse))) , mux_105_cse},
      (else_7_if_div_9cyc_st_7[1]) | (else_7_if_div_9cyc_st_7[0]) | if_7_equal_svs_st_7
      | (~ main_stage_0_8) | (else_7_if_div_9cyc_st_7[2]) | (else_7_if_div_9cyc_st_7[3]));
  assign mux_122_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_46))) , and_tmp_46},
      or_tmp_184);
  assign and_3312_cse = (mux_122_nl) & and_dcpl_3158 & and_dcpl_3249 & (~ (else_7_if_div_9cyc_st_2[2]));
  assign mux_123_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_47))) , and_tmp_47},
      or_tmp_184);
  assign and_3320_cse = or_tmp_15 & (mux_123_nl) & and_dcpl_3258 & and_dcpl_3162;
  assign and_3329_cse = or_tmp_23 & or_831_cse & or_833_cse & mux_124_cse & and_dcpl_3264
      & and_dcpl_3168;
  assign and_3339_cse = or_tmp_33 & ((~ or_tmp_34) | (else_7_if_div_9cyc_st_4[3])
      | (else_7_if_div_9cyc_st_4[2]) | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0]))
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_831_cse & or_833_cse & mux_124_cse
      & and_dcpl_3270 & and_dcpl_3174;
  assign mux_129_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_60))) , and_tmp_60},
      or_835_cse);
  assign and_3361_cse = ((~ or_tmp_60) | (else_7_if_div_9cyc_st_6[3]) | (else_7_if_div_9cyc_st_6[2])
      | (else_7_if_div_9cyc_st_6[1]) | (~ (else_7_if_div_9cyc_st_6[0])) | (~ main_stage_0_7)
      | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (else_7_if_div_9cyc_st_5[3]) | (else_7_if_div_9cyc_st_5[2])
      | (else_7_if_div_9cyc_st_5[1]) | (~ (else_7_if_div_9cyc_st_5[0])) | (~ main_stage_0_6)
      | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0])) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_831_cse & or_833_cse & (mux_129_nl) & and_dcpl_3188
      & and_dcpl_3280;
  assign mux_127_nl = MUX_s_1_2_2({and_3347_cse , (~(or_tmp_58 | (~ and_3347_cse)))},
      main_stage_0_6);
  assign mux_128_nl = MUX_s_1_2_2({(mux_127_nl) , and_3347_cse}, or_tmp_221);
  assign and_3349_cse = or_tmp_45 & (mux_128_nl) & and_dcpl_3276 & and_dcpl_3180;
  assign mux_135_cse = MUX_s_1_2_2({(~(or_tmp_94 | (~ mux_134_cse))) , mux_134_cse},
      (else_7_if_div_9cyc_st_7[1]) | (~ (else_7_if_div_9cyc_st_7[0])) | if_7_equal_svs_st_7
      | (~ main_stage_0_8) | (else_7_if_div_9cyc_st_7[2]) | (else_7_if_div_9cyc_st_7[3]));
  assign mux_151_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_92))) , and_tmp_92},
      or_tmp_359);
  assign and_3452_cse = (mux_151_nl) & and_dcpl_3158 & and_dcpl_3343 & (~ (else_7_if_div_9cyc_st_2[2]));
  assign mux_152_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_93))) , and_tmp_93},
      or_tmp_359);
  assign and_3460_cse = or_tmp_15 & (mux_152_nl) & and_dcpl_3164 & and_dcpl_3350;
  assign and_3469_cse = or_tmp_23 & or_1036_cse & or_1038_cse & mux_153_cse & and_dcpl_3170
      & and_dcpl_3356;
  assign and_3479_cse = or_tmp_33 & ((~ or_tmp_34) | (else_7_if_div_9cyc_st_4[3])
      | (else_7_if_div_9cyc_st_4[2]) | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1036_cse & or_1038_cse & mux_153_cse
      & and_dcpl_3176 & and_dcpl_3362;
  assign mux_158_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_106))) , and_tmp_106},
      or_1040_cse);
  assign and_3501_cse = ((~ or_tmp_60) | (else_7_if_div_9cyc_st_6[3]) | (else_7_if_div_9cyc_st_6[2])
      | (~ (else_7_if_div_9cyc_st_6[1])) | (else_7_if_div_9cyc_st_6[0]) | (~ main_stage_0_7)
      | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (else_7_if_div_9cyc_st_5[3]) | (else_7_if_div_9cyc_st_5[2])
      | (~ (else_7_if_div_9cyc_st_5[1])) | (else_7_if_div_9cyc_st_5[0]) | (~ main_stage_0_6)
      | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (else_7_if_div_9cyc_st_4[3]) | (else_7_if_div_9cyc_st_4[2])
      | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0]) | (~ main_stage_0_5)
      | if_7_equal_svs_st_4) & or_1036_cse & or_1038_cse & (mux_158_nl) & and_dcpl_3188
      & and_dcpl_3374;
  assign mux_156_nl = MUX_s_1_2_2({and_3487_cse , (~(or_tmp_58 | (~ and_3487_cse)))},
      main_stage_0_6);
  assign mux_157_nl = MUX_s_1_2_2({(mux_156_nl) , and_3487_cse}, or_tmp_396);
  assign and_3489_cse = or_tmp_45 & (mux_157_nl) & and_dcpl_3182 & and_dcpl_3368;
  assign mux_164_cse = MUX_s_1_2_2({(~(or_tmp_94 | (~ mux_163_cse))) , mux_163_cse},
      (~ (else_7_if_div_9cyc_st_7[1])) | (else_7_if_div_9cyc_st_7[0]) | if_7_equal_svs_st_7
      | (~ main_stage_0_8) | (else_7_if_div_9cyc_st_7[2]) | (else_7_if_div_9cyc_st_7[3]));
  assign mux_180_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_138))) , and_tmp_138},
      or_tmp_534);
  assign and_3592_cse = (mux_180_nl) & and_dcpl_3158 & and_dcpl_3437 & (~ (else_7_if_div_9cyc_st_2[2]));
  assign mux_181_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_139))) , and_tmp_139},
      or_tmp_534);
  assign and_3600_cse = or_tmp_15 & (mux_181_nl) & and_dcpl_3258 & and_dcpl_3350;
  assign and_3609_cse = or_tmp_23 & or_1241_cse & or_1243_cse & mux_182_cse & and_dcpl_3264
      & and_dcpl_3356;
  assign and_3619_cse = or_tmp_33 & ((~ or_tmp_34) | (else_7_if_div_9cyc_st_4[3])
      | (else_7_if_div_9cyc_st_4[2]) | (~ (else_7_if_div_9cyc_st_4[1])) | (~ (else_7_if_div_9cyc_st_4[0]))
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1241_cse & or_1243_cse & mux_182_cse
      & and_dcpl_3270 & and_dcpl_3362;
  assign mux_187_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_152))) , and_tmp_152},
      or_1245_cse);
  assign and_3641_cse = ((~ or_tmp_60) | (else_7_if_div_9cyc_st_6[3]) | (else_7_if_div_9cyc_st_6[2])
      | (~ (else_7_if_div_9cyc_st_6[1])) | (~ (else_7_if_div_9cyc_st_6[0])) | (~
      main_stage_0_7) | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (else_7_if_div_9cyc_st_5[3])
      | (else_7_if_div_9cyc_st_5[2]) | (~ (else_7_if_div_9cyc_st_5[1])) | (~ (else_7_if_div_9cyc_st_5[0]))
      | (~ main_stage_0_6) | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (else_7_if_div_9cyc_st_4[3])
      | (else_7_if_div_9cyc_st_4[2]) | (~ (else_7_if_div_9cyc_st_4[1])) | (~ (else_7_if_div_9cyc_st_4[0]))
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1241_cse & or_1243_cse & (mux_187_nl)
      & and_dcpl_3188 & and_dcpl_3468;
  assign mux_185_nl = MUX_s_1_2_2({and_3627_cse , (~(or_tmp_58 | (~ and_3627_cse)))},
      main_stage_0_6);
  assign mux_186_nl = MUX_s_1_2_2({(mux_185_nl) , and_3627_cse}, or_tmp_571);
  assign and_3629_cse = or_tmp_45 & (mux_186_nl) & and_dcpl_3276 & and_dcpl_3368;
  assign mux_193_nl = MUX_s_1_2_2({mux_192_cse , (~(or_tmp_94 | (~ mux_192_cse)))},
      main_stage_0_8);
  assign mux_194_cse = MUX_s_1_2_2({(mux_193_nl) , mux_192_cse}, (else_7_if_div_9cyc_st_7[3])
      | (else_7_if_div_9cyc_st_7[2]) | (~ (else_7_if_div_9cyc_st_7[1])) | (~ (else_7_if_div_9cyc_st_7[0]))
      | if_7_equal_svs_st_7);
  assign mux_211_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_184))) , and_tmp_184},
      or_tmp_709);
  assign and_3732_cse = (mux_211_nl) & and_dcpl_3158 & and_dcpl_3155 & (else_7_if_div_9cyc_st_2[2]);
  assign mux_212_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_185))) , and_tmp_185},
      or_tmp_709);
  assign and_3740_cse = or_tmp_15 & (mux_212_nl) & and_dcpl_3164 & and_dcpl_3538;
  assign and_3749_cse = or_tmp_23 & or_1446_cse & or_1448_cse & mux_213_cse & and_dcpl_3170
      & and_dcpl_3544;
  assign and_3759_cse = or_tmp_33 & ((~ or_tmp_34) | (else_7_if_div_9cyc_st_4[3])
      | (~ (else_7_if_div_9cyc_st_4[2])) | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1446_cse & or_1448_cse & mux_213_cse
      & and_dcpl_3176 & and_dcpl_3550;
  assign mux_218_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_198))) , and_tmp_198},
      or_1450_cse);
  assign and_3781_cse = ((~ or_tmp_60) | (else_7_if_div_9cyc_st_6[3]) | (~ (else_7_if_div_9cyc_st_6[2]))
      | (else_7_if_div_9cyc_st_6[1]) | (else_7_if_div_9cyc_st_6[0]) | (~ main_stage_0_7)
      | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (else_7_if_div_9cyc_st_5[3]) | (~
      (else_7_if_div_9cyc_st_5[2])) | (else_7_if_div_9cyc_st_5[1]) | (else_7_if_div_9cyc_st_5[0])
      | (~ main_stage_0_6) | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (else_7_if_div_9cyc_st_4[3])
      | (~ (else_7_if_div_9cyc_st_4[2])) | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1446_cse & or_1448_cse & (mux_218_nl)
      & and_dcpl_3564 & and_dcpl_3186;
  assign mux_216_nl = MUX_s_1_2_2({and_3767_cse , (~(or_tmp_58 | (~ and_3767_cse)))},
      main_stage_0_6);
  assign mux_217_nl = MUX_s_1_2_2({(mux_216_nl) , and_3767_cse}, or_tmp_746);
  assign and_3769_cse = or_tmp_45 & (mux_217_nl) & and_dcpl_3182 & and_dcpl_3556;
  assign mux_224_cse = MUX_s_1_2_2({(~(or_tmp_94 | (~ mux_223_cse))) , mux_223_cse},
      (else_7_if_div_9cyc_st_7[1]) | (else_7_if_div_9cyc_st_7[0]) | if_7_equal_svs_st_7
      | (~ main_stage_0_8) | (~ (else_7_if_div_9cyc_st_7[2])) | (else_7_if_div_9cyc_st_7[3]));
  assign mux_240_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_230))) , and_tmp_230},
      or_tmp_884);
  assign and_3872_cse = (mux_240_nl) & and_dcpl_3158 & and_dcpl_3249 & (else_7_if_div_9cyc_st_2[2]);
  assign mux_241_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_231))) , and_tmp_231},
      or_tmp_884);
  assign and_3880_cse = or_tmp_15 & (mux_241_nl) & and_dcpl_3258 & and_dcpl_3538;
  assign and_3889_cse = or_tmp_23 & or_1651_cse & or_1653_cse & mux_242_cse & and_dcpl_3264
      & and_dcpl_3544;
  assign and_3899_cse = or_tmp_33 & ((~ or_tmp_34) | (else_7_if_div_9cyc_st_4[3])
      | (~ (else_7_if_div_9cyc_st_4[2])) | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0]))
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1651_cse & or_1653_cse & mux_242_cse
      & and_dcpl_3270 & and_dcpl_3550;
  assign mux_247_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_244))) , and_tmp_244},
      or_1655_cse);
  assign and_3921_cse = ((~ or_tmp_60) | (else_7_if_div_9cyc_st_6[3]) | (~ (else_7_if_div_9cyc_st_6[2]))
      | (else_7_if_div_9cyc_st_6[1]) | (~ (else_7_if_div_9cyc_st_6[0])) | (~ main_stage_0_7)
      | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (else_7_if_div_9cyc_st_5[3]) | (~
      (else_7_if_div_9cyc_st_5[2])) | (else_7_if_div_9cyc_st_5[1]) | (~ (else_7_if_div_9cyc_st_5[0]))
      | (~ main_stage_0_6) | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (else_7_if_div_9cyc_st_4[3])
      | (~ (else_7_if_div_9cyc_st_4[2])) | (else_7_if_div_9cyc_st_4[1]) | (~ (else_7_if_div_9cyc_st_4[0]))
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1651_cse & or_1653_cse & (mux_247_nl)
      & and_dcpl_3564 & and_dcpl_3280;
  assign mux_245_nl = MUX_s_1_2_2({and_3907_cse , (~(or_tmp_58 | (~ and_3907_cse)))},
      main_stage_0_6);
  assign mux_246_nl = MUX_s_1_2_2({(mux_245_nl) , and_3907_cse}, or_tmp_921);
  assign and_3909_cse = or_tmp_45 & (mux_246_nl) & and_dcpl_3276 & and_dcpl_3556;
  assign mux_253_cse = MUX_s_1_2_2({(~(or_tmp_94 | (~ mux_252_cse))) , mux_252_cse},
      (else_7_if_div_9cyc_st_7[1]) | (~ (else_7_if_div_9cyc_st_7[0])) | if_7_equal_svs_st_7
      | (~ main_stage_0_8) | (~ (else_7_if_div_9cyc_st_7[2])) | (else_7_if_div_9cyc_st_7[3]));
  assign mux_269_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_276))) , and_tmp_276},
      or_tmp_1059);
  assign and_4012_cse = (mux_269_nl) & and_dcpl_3158 & and_dcpl_3343 & (else_7_if_div_9cyc_st_2[2]);
  assign mux_270_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_277))) , and_tmp_277},
      or_tmp_1059);
  assign and_4020_cse = or_tmp_15 & (mux_270_nl) & and_dcpl_3164 & and_dcpl_3726;
  assign and_4029_cse = or_tmp_23 & or_1856_cse & or_1858_cse & mux_271_cse & and_dcpl_3170
      & and_dcpl_3732;
  assign and_4039_cse = or_tmp_33 & ((~ or_tmp_34) | (else_7_if_div_9cyc_st_4[3])
      | (~ (else_7_if_div_9cyc_st_4[2])) | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1856_cse & or_1858_cse & mux_271_cse
      & and_dcpl_3176 & and_dcpl_3738;
  assign mux_276_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_290))) , and_tmp_290},
      or_1860_cse);
  assign and_4061_cse = ((~ or_tmp_60) | (else_7_if_div_9cyc_st_6[3]) | (~ (else_7_if_div_9cyc_st_6[2]))
      | (~ (else_7_if_div_9cyc_st_6[1])) | (else_7_if_div_9cyc_st_6[0]) | (~ main_stage_0_7)
      | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (else_7_if_div_9cyc_st_5[3]) | (~
      (else_7_if_div_9cyc_st_5[2])) | (~ (else_7_if_div_9cyc_st_5[1])) | (else_7_if_div_9cyc_st_5[0])
      | (~ main_stage_0_6) | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (else_7_if_div_9cyc_st_4[3])
      | (~ (else_7_if_div_9cyc_st_4[2])) | (~ (else_7_if_div_9cyc_st_4[1])) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_1856_cse & or_1858_cse & (mux_276_nl)
      & and_dcpl_3564 & and_dcpl_3374;
  assign mux_274_nl = MUX_s_1_2_2({and_4047_cse , (~(or_tmp_58 | (~ and_4047_cse)))},
      main_stage_0_6);
  assign mux_275_nl = MUX_s_1_2_2({(mux_274_nl) , and_4047_cse}, or_tmp_1096);
  assign and_4049_cse = or_tmp_45 & (mux_275_nl) & and_dcpl_3182 & and_dcpl_3744;
  assign mux_282_cse = MUX_s_1_2_2({(~(or_tmp_94 | (~ mux_281_cse))) , mux_281_cse},
      (~ (else_7_if_div_9cyc_st_7[1])) | (else_7_if_div_9cyc_st_7[0]) | if_7_equal_svs_st_7
      | (~ main_stage_0_8) | (~ (else_7_if_div_9cyc_st_7[2])) | (else_7_if_div_9cyc_st_7[3]));
  assign mux_298_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_322))) , and_tmp_322},
      or_tmp_1234);
  assign and_4152_cse = (mux_298_nl) & and_dcpl_3158 & and_dcpl_3437 & (else_7_if_div_9cyc_st_2[2]);
  assign mux_299_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ and_tmp_323))) , and_tmp_323},
      or_tmp_1234);
  assign and_4160_cse = or_tmp_15 & (mux_299_nl) & and_dcpl_3258 & and_dcpl_3726;
  assign and_4169_cse = or_tmp_23 & or_2061_cse & nand_33_cse & mux_302_cse & and_dcpl_3264
      & and_dcpl_3732;
  assign and_4179_cse = or_tmp_33 & (~(or_tmp_34 & (~ (else_7_if_div_9cyc_st_4[3]))
      & (else_7_if_div_9cyc_st_4[2]) & (else_7_if_div_9cyc_st_4[1]) & (else_7_if_div_9cyc_st_4[0])
      & main_stage_0_5 & (~ if_7_equal_svs_st_4))) & or_2061_cse & nand_33_cse &
      mux_302_cse & and_dcpl_3270 & and_dcpl_3738;
  assign mux_305_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_4195_cse))) , and_4195_cse},
      or_2065_cse);
  assign and_4201_cse = (~(or_tmp_60 & (~ (else_7_if_div_9cyc_st_6[3])) & (else_7_if_div_9cyc_st_6[2])
      & (else_7_if_div_9cyc_st_6[1]) & (else_7_if_div_9cyc_st_6[0]) & main_stage_0_7
      & (~ if_7_equal_svs_st_6))) & (~(or_tmp_33 & (~ (else_7_if_div_9cyc_st_5[3]))
      & (else_7_if_div_9cyc_st_5[2]) & (else_7_if_div_9cyc_st_5[1]) & (else_7_if_div_9cyc_st_5[0])
      & main_stage_0_6 & (~ if_7_equal_svs_st_5))) & (~(or_tmp_64 & (~ (else_7_if_div_9cyc_st_4[3]))
      & (else_7_if_div_9cyc_st_4[2]) & (else_7_if_div_9cyc_st_4[1]) & (else_7_if_div_9cyc_st_4[0])
      & main_stage_0_5 & (~ if_7_equal_svs_st_4))) & or_2061_cse & nand_33_cse &
      (mux_305_nl) & and_dcpl_3564 & and_dcpl_3468;
  assign mux_303_nl = MUX_s_1_2_2({and_4187_cse , (~(or_tmp_58 | (~ and_4187_cse)))},
      main_stage_0_6);
  assign mux_304_nl = MUX_s_1_2_2({(mux_303_nl) , and_4187_cse}, or_tmp_1271);
  assign and_4189_cse = or_tmp_45 & (mux_304_nl) & and_dcpl_3276 & and_dcpl_3744;
  assign mux_311_nl = MUX_s_1_2_2({mux_310_cse , (~(or_tmp_94 | (~ mux_310_cse)))},
      main_stage_0_8);
  assign mux_312_cse = MUX_s_1_2_2({(mux_311_nl) , mux_310_cse}, (else_7_if_div_9cyc_st_7[3])
      | (~ (else_7_if_div_9cyc_st_7[2])) | (~ (else_7_if_div_9cyc_st_7[1])) | (~
      (else_7_if_div_9cyc_st_7[0])) | if_7_equal_svs_st_7);
  assign mux_330_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ mux_tmp_246))) , mux_tmp_246},
      or_tmp_1409);
  assign and_4291_cse = (mux_330_nl) & and_1994_cse & (else_7_if_div_9cyc_st_2[3])
      & and_dcpl_3156;
  assign mux_332_nl = MUX_s_1_2_2({(~(or_tmp_7 | (~ mux_tmp_248))) , mux_tmp_248},
      or_tmp_1409);
  assign and_4298_cse = or_tmp_15 & (mux_332_nl) & and_dcpl_3164 & and_dcpl_3161
      & (else_7_if_div_9cyc_st_3[3]);
  assign and_4307_cse = or_tmp_23 & or_2269_cse & or_2271_cse & mux_333_cse & and_dcpl_3170
      & and_dcpl_3167 & (else_7_if_div_9cyc_st_4[3]);
  assign and_4317_cse = or_tmp_33 & ((~ or_tmp_34) | (~ (else_7_if_div_9cyc_st_4[3]))
      | (else_7_if_div_9cyc_st_4[2]) | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_2269_cse & or_2271_cse & mux_333_cse
      & and_dcpl_3176 & and_dcpl_3173 & (else_7_if_div_9cyc_st_5[3]);
  assign mux_338_nl = MUX_s_1_2_2({(~(main_stage_0_3 | (~ and_tmp_380))) , and_tmp_380},
      or_2273_cse);
  assign and_4339_cse = ((~ or_tmp_60) | (~ (else_7_if_div_9cyc_st_6[3])) | (else_7_if_div_9cyc_st_6[2])
      | (else_7_if_div_9cyc_st_6[1]) | (else_7_if_div_9cyc_st_6[0]) | (~ main_stage_0_7)
      | if_7_equal_svs_st_6) & ((~ or_tmp_33) | (~ (else_7_if_div_9cyc_st_5[3]))
      | (else_7_if_div_9cyc_st_5[2]) | (else_7_if_div_9cyc_st_5[1]) | (else_7_if_div_9cyc_st_5[0])
      | (~ main_stage_0_6) | if_7_equal_svs_st_5) & ((~ or_tmp_64) | (~ (else_7_if_div_9cyc_st_4[3]))
      | (else_7_if_div_9cyc_st_4[2]) | (else_7_if_div_9cyc_st_4[1]) | (else_7_if_div_9cyc_st_4[0])
      | (~ main_stage_0_5) | if_7_equal_svs_st_4) & or_2269_cse & or_2271_cse & (mux_338_nl)
      & and_dcpl_3188 & (else_7_if_div_9cyc_st_7[3]) & (~ (else_7_if_div_9cyc_st_7[0]))
      & (~ (else_7_if_div_9cyc_st_7[1]));
  assign mux_336_nl = MUX_s_1_2_2({and_4325_cse , (~(or_tmp_58 | (~ and_4325_cse)))},
      main_stage_0_6);
  assign mux_337_nl = MUX_s_1_2_2({(mux_336_nl) , and_4325_cse}, or_tmp_1449);
  assign and_4327_cse = or_tmp_45 & (mux_337_nl) & and_dcpl_3182 & and_dcpl_3179
      & (else_7_if_div_9cyc_st_6[3]);
  assign mux_344_nl = MUX_s_1_2_2({mux_343_cse , (~(or_tmp_94 | (~ mux_343_cse)))},
      else_7_if_div_9cyc_st_7[3]);
  assign mux_345_cse = MUX_s_1_2_2({(mux_344_nl) , mux_343_cse}, (else_7_if_div_9cyc_st_7[1])
      | (else_7_if_div_9cyc_st_7[0]) | if_7_equal_svs_st_7 | (~ main_stage_0_8) |
      (else_7_if_div_9cyc_st_7[2]));
  assign and_5652_cse = mux_466_cse & and_dcpl_4020 & (else_7_if_1_div_9cyc_st_4[3])
      & (~ (else_7_if_1_div_9cyc_st_4[0])) & (~ (else_7_if_1_div_9cyc_st_4[1]));
  assign and_5659_cse = mux_471_cse & and_878_cse & else_7_equal_svs_st_5 & (else_7_if_1_div_9cyc_st_5[3])
      & and_dcpl_4024;
  assign mux_472_nl = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_5[3]) | (~ mux_471_cse)))
      , mux_471_cse}, or_tmp_2252);
  assign and_5666_cse = (mux_472_nl) & and_dcpl_4034 & (else_7_if_1_div_9cyc_st_6[3])
      & (~ (else_7_if_1_div_9cyc_st_6[0])) & (~ (else_7_if_1_div_9cyc_st_6[1]));
  assign and_5674_cse = mux_482_cse & and_dcpl_4041 & (else_7_if_1_div_9cyc_st_7[3])
      & (~ (else_7_if_1_div_9cyc_st_7[0])) & (~ (else_7_if_1_div_9cyc_st_7[1]));
  assign mux_483_cse = MUX_s_1_2_2({(~((else_7_if_1_div_9cyc_st_7[3]) | (~ mux_482_cse)))
      , mux_482_cse}, (~ main_stage_0_8) | if_7_equal_svs_st_7 | (~ else_7_equal_svs_st_7)
      | (else_7_if_1_div_9cyc_st_7[0]) | (else_7_if_1_div_9cyc_st_7[1]) | (else_7_if_1_div_9cyc_st_7[2]));
  assign mux_607_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ mux_tmp_523)))
      , mux_tmp_523}, or_tmp_2993);
  assign and_7108_cse = (mux_607_nl) & and_dcpl_4997 & (~ (else_7_else_1_if_div_9cyc_st_4[2]))
      & (else_7_else_1_if_div_9cyc_st_4[3]) & and_dcpl_1350;
  assign mux_611_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ mux_610_cse)))
      , mux_610_cse}, or_tmp_2993);
  assign and_7116_cse = (mux_611_nl) & and_dcpl_5005 & (~ (else_7_else_1_if_div_9cyc_st_5[2]))
      & (else_7_else_1_if_div_9cyc_st_5[3]) & and_dcpl_978;
  assign mux_616_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ mux_615_cse)))
      , mux_615_cse}, or_tmp_2993);
  assign and_7124_cse = (mux_616_nl) & and_dcpl_5013 & (~ (else_7_else_1_if_div_9cyc_st_6[2]))
      & (else_7_else_1_if_div_9cyc_st_6[3]) & and_dcpl_606;
  assign mux_622_nl = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ mux_621_cse)))
      , mux_621_cse}, or_tmp_2993);
  assign and_7132_cse = (mux_622_nl) & and_dcpl_5021 & (~ (else_7_else_1_if_div_9cyc_st_7[2]))
      & (else_7_else_1_if_div_9cyc_st_7[3]) & and_dcpl_234;
  assign mux_628_cse = MUX_s_1_2_2({(~(else_7_else_1_equal_svs_1 | (~ mux_627_cse)))
      , mux_627_cse}, or_tmp_2993);
  assign and_8682_cse = or_tmp_3659 & mux_659_cse & and_1246_cse & (~ (else_7_else_1_else_div_9cyc_st_5[2]))
      & (else_7_else_1_else_div_9cyc_st_5[3]) & and_dcpl_1107;
  assign and_8691_cse = or_tmp_3659 & mux_664_cse & and_874_cse & (~ (else_7_else_1_else_div_9cyc_st_6[2]))
      & (else_7_else_1_else_div_9cyc_st_6[3]) & and_dcpl_735;
  assign mux_665_nl = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_6[3]) | (~
      mux_664_cse))) , mux_664_cse}, or_tmp_3688);
  assign and_8700_cse = or_tmp_3659 & (mux_665_nl) & and_502_cse & (~ (else_7_else_1_else_div_9cyc_st_7[2]))
      & (else_7_else_1_else_div_9cyc_st_7[3]) & and_dcpl_363;
  assign mux_670_nl = MUX_s_1_2_2({(~((else_7_else_1_else_div_9cyc_st_7[3]) | (~
      and_8701_cse))) , and_8701_cse}, (~ main_stage_0_8) | if_7_equal_svs_st_7 |
      else_7_equal_svs_st_7 | else_7_else_1_equal_svs_st_7 | (else_7_else_1_else_div_9cyc_st_7[0])
      | (else_7_else_1_else_div_9cyc_st_7[1]) | (else_7_else_1_else_div_9cyc_st_7[2]));
  assign and_8702_cse = or_tmp_3659 & (mux_670_nl);
  always @(posedge clk) begin
    if ( rst ) begin
      V_OUT_rsc_mgc_out_stdreg_d <= 32'b0;
      S_OUT_rsc_mgc_out_stdreg_d <= 32'b0;
      H_OUT_rsc_mgc_out_stdreg_d <= 32'b0;
      else_7_acc_2_psp_sg1_sva <= 16'b0;
      else_7_if_div_tmp_duc_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_9 <= 4'b0;
      h_2_sva_duc <= 30'b0;
      else_7_if_1_div_9cyc_st_9 <= 4'b0;
      div_sdt_2_sva_duc <= 30'b0;
      div_sdt_3_sva_duc <= 30'b0;
      else_7_else_1_if_div_9cyc_st_9 <= 4'b0;
      else_7_else_1_else_div_9cyc_st_9 <= 4'b0;
      else_7_else_1_equal_svs_st_9 <= 1'b0;
      else_7_and_5_itm_9 <= 1'b0;
      else_7_equal_svs_9 <= 1'b0;
      unequal_tmp_9 <= 1'b0;
      max_sg1_lpi_dfm_3_st_9 <= 16'b0;
      slc_3_itm_9 <= 15'b0;
      if_7_equal_svs_9 <= 1'b0;
      max_conc_4_tmp_mut_24_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_24_sg1 <= 16'b0;
      max_conc_4_tmp_mut_32_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_32_sg1 <= 16'b0;
      max_conc_4_tmp_mut_40_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_40_sg1 <= 16'b0;
      max_conc_4_tmp_mut_48_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_48_sg1 <= 16'b0;
      max_conc_4_tmp_mut_56_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_56_sg1 <= 16'b0;
      max_conc_4_tmp_mut_64_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_64_sg1 <= 16'b0;
      max_conc_4_tmp_mut_72_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_72_sg1 <= 16'b0;
      max_conc_4_tmp_mut_80_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_80_sg1 <= 16'b0;
      max_conc_4_tmp_mut_16_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_16_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_8 <= 4'b0;
      delta_conc_1_tmp_mut_24_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_24_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_32_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_32_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_40_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_40_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_48_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_48_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_56_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_56_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_64_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_64_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_72_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_72_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_80_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_80_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_16_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_16_sg1 <= 17'b0;
      else_7_if_1_div_9cyc_st_8 <= 4'b0;
      delta_conc_2_tmp_mut_16_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_16_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_24_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_24_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_32_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_32_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_40_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_40_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_48_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_48_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_56_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_56_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_64_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_64_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_72_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_72_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_80_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_80_sg1 <= 17'b0;
      else_7_else_1_if_div_9cyc_st_8 <= 4'b0;
      delta_conc_3_tmp_mut_16_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_16_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_24_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_24_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_32_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_32_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_40_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_40_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_48_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_48_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_56_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_56_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_64_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_64_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_72_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_72_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_80_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_80_sg1 <= 17'b0;
      else_7_else_1_else_div_9cyc_st_8 <= 4'b0;
      else_7_else_1_equal_svs_st_8 <= 1'b0;
      else_7_equal_svs_st_8 <= 1'b0;
      max_sg1_lpi_dfm_3_st_8 <= 16'b0;
      if_7_equal_svs_st_8 <= 1'b0;
      max_conc_4_tmp_mut_23_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_23_sg1 <= 16'b0;
      max_conc_4_tmp_mut_31_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_31_sg1 <= 16'b0;
      max_conc_4_tmp_mut_39_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_39_sg1 <= 16'b0;
      max_conc_4_tmp_mut_47_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_47_sg1 <= 16'b0;
      max_conc_4_tmp_mut_55_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_55_sg1 <= 16'b0;
      max_conc_4_tmp_mut_63_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_63_sg1 <= 16'b0;
      max_conc_4_tmp_mut_71_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_71_sg1 <= 16'b0;
      max_conc_4_tmp_mut_79_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_79_sg1 <= 16'b0;
      max_conc_4_tmp_mut_15_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_15_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_7 <= 4'b0;
      delta_conc_1_tmp_mut_23_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_23_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_31_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_31_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_39_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_39_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_47_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_47_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_55_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_55_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_63_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_63_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_71_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_71_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_79_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_79_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_15_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_15_sg1 <= 17'b0;
      else_7_if_1_div_9cyc_st_7 <= 4'b0;
      delta_conc_2_tmp_mut_15_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_15_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_23_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_23_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_31_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_31_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_39_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_39_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_47_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_47_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_55_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_55_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_63_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_63_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_71_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_71_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_79_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_79_sg1 <= 17'b0;
      else_7_else_1_if_div_9cyc_st_7 <= 4'b0;
      delta_conc_3_tmp_mut_15_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_15_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_23_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_23_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_31_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_31_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_39_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_39_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_47_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_47_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_55_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_55_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_63_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_63_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_71_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_71_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_79_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_79_sg1 <= 17'b0;
      else_7_else_1_else_div_9cyc_st_7 <= 4'b0;
      else_7_else_1_equal_svs_st_7 <= 1'b0;
      else_7_equal_svs_st_7 <= 1'b0;
      max_sg1_lpi_dfm_3_st_7 <= 16'b0;
      if_7_equal_svs_st_7 <= 1'b0;
      max_conc_4_tmp_mut_22_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_22_sg1 <= 16'b0;
      max_conc_4_tmp_mut_30_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_30_sg1 <= 16'b0;
      max_conc_4_tmp_mut_38_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_38_sg1 <= 16'b0;
      max_conc_4_tmp_mut_46_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_46_sg1 <= 16'b0;
      max_conc_4_tmp_mut_54_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_54_sg1 <= 16'b0;
      max_conc_4_tmp_mut_62_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_62_sg1 <= 16'b0;
      max_conc_4_tmp_mut_70_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_70_sg1 <= 16'b0;
      max_conc_4_tmp_mut_78_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_78_sg1 <= 16'b0;
      max_conc_4_tmp_mut_14_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_14_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_6 <= 4'b0;
      delta_conc_1_tmp_mut_22_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_22_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_30_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_30_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_38_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_38_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_46_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_46_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_54_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_54_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_62_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_62_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_70_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_70_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_78_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_78_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_14_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_14_sg1 <= 17'b0;
      else_7_if_1_div_9cyc_st_6 <= 4'b0;
      delta_conc_2_tmp_mut_14_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_14_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_22_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_22_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_30_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_30_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_38_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_38_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_46_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_46_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_54_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_54_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_62_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_62_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_70_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_70_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_78_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_78_sg1 <= 17'b0;
      else_7_else_1_if_div_9cyc_st_6 <= 4'b0;
      delta_conc_3_tmp_mut_14_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_14_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_22_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_22_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_30_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_30_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_38_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_38_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_46_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_46_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_54_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_54_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_62_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_62_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_70_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_70_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_78_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_78_sg1 <= 17'b0;
      else_7_else_1_else_div_9cyc_st_6 <= 4'b0;
      else_7_else_1_equal_svs_st_6 <= 1'b0;
      else_7_equal_svs_st_6 <= 1'b0;
      max_sg1_lpi_dfm_3_st_6 <= 16'b0;
      if_7_equal_svs_st_6 <= 1'b0;
      max_conc_4_tmp_mut_21_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_21_sg1 <= 16'b0;
      max_conc_4_tmp_mut_29_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_29_sg1 <= 16'b0;
      max_conc_4_tmp_mut_37_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_37_sg1 <= 16'b0;
      max_conc_4_tmp_mut_45_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_45_sg1 <= 16'b0;
      max_conc_4_tmp_mut_53_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_53_sg1 <= 16'b0;
      max_conc_4_tmp_mut_61_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_61_sg1 <= 16'b0;
      max_conc_4_tmp_mut_69_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_69_sg1 <= 16'b0;
      max_conc_4_tmp_mut_77_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_77_sg1 <= 16'b0;
      max_conc_4_tmp_mut_13_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_13_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_5 <= 4'b0;
      delta_conc_1_tmp_mut_21_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_21_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_29_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_29_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_37_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_37_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_45_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_45_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_53_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_53_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_61_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_61_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_69_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_69_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_77_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_77_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_13_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_13_sg1 <= 17'b0;
      else_7_if_1_div_9cyc_st_5 <= 4'b0;
      delta_conc_2_tmp_mut_13_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_13_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_21_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_21_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_29_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_29_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_37_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_37_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_45_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_45_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_53_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_53_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_61_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_61_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_69_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_69_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_77_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_77_sg1 <= 17'b0;
      else_7_else_1_if_div_9cyc_st_5 <= 4'b0;
      delta_conc_3_tmp_mut_13_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_13_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_21_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_21_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_29_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_29_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_37_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_37_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_45_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_45_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_53_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_53_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_61_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_61_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_69_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_69_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_77_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_77_sg1 <= 17'b0;
      else_7_else_1_else_div_9cyc_st_5 <= 4'b0;
      else_7_else_1_equal_svs_st_5 <= 1'b0;
      else_7_equal_svs_st_5 <= 1'b0;
      max_sg1_lpi_dfm_3_st_5 <= 16'b0;
      if_7_equal_svs_st_5 <= 1'b0;
      max_conc_4_tmp_mut_20_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_20_sg1 <= 16'b0;
      max_conc_4_tmp_mut_28_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_28_sg1 <= 16'b0;
      max_conc_4_tmp_mut_36_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_36_sg1 <= 16'b0;
      max_conc_4_tmp_mut_44_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_44_sg1 <= 16'b0;
      max_conc_4_tmp_mut_52_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_52_sg1 <= 16'b0;
      max_conc_4_tmp_mut_60_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_60_sg1 <= 16'b0;
      max_conc_4_tmp_mut_68_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_68_sg1 <= 16'b0;
      max_conc_4_tmp_mut_76_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_76_sg1 <= 16'b0;
      max_conc_4_tmp_mut_12_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_12_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_4 <= 4'b0;
      delta_conc_1_tmp_mut_20_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_20_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_28_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_28_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_36_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_36_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_44_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_44_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_52_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_52_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_60_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_60_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_68_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_68_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_76_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_76_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_12_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_12_sg1 <= 17'b0;
      else_7_if_1_div_9cyc_st_4 <= 4'b0;
      delta_conc_2_tmp_mut_12_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_12_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_20_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_20_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_28_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_28_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_36_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_36_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_44_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_44_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_52_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_52_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_60_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_60_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_68_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_68_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_76_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_76_sg1 <= 17'b0;
      else_7_else_1_if_div_9cyc_st_4 <= 4'b0;
      delta_conc_3_tmp_mut_12_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_12_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_20_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_20_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_28_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_28_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_36_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_36_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_44_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_44_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_52_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_52_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_60_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_60_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_68_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_68_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_76_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_76_sg1 <= 17'b0;
      else_7_else_1_else_div_9cyc_st_4 <= 4'b0;
      else_7_else_1_equal_svs_st_4 <= 1'b0;
      else_7_equal_svs_st_4 <= 1'b0;
      max_sg1_lpi_dfm_3_st_4 <= 16'b0;
      if_7_equal_svs_st_4 <= 1'b0;
      max_conc_4_tmp_mut_19_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_19_sg1 <= 16'b0;
      max_conc_4_tmp_mut_27_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_27_sg1 <= 16'b0;
      max_conc_4_tmp_mut_35_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_35_sg1 <= 16'b0;
      max_conc_4_tmp_mut_43_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_43_sg1 <= 16'b0;
      max_conc_4_tmp_mut_51_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_51_sg1 <= 16'b0;
      max_conc_4_tmp_mut_59_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_59_sg1 <= 16'b0;
      max_conc_4_tmp_mut_67_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_67_sg1 <= 16'b0;
      max_conc_4_tmp_mut_75_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_75_sg1 <= 16'b0;
      max_conc_4_tmp_mut_11_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_11_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_3 <= 4'b0;
      delta_conc_1_tmp_mut_19_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_19_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_27_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_27_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_35_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_35_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_43_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_43_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_51_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_51_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_59_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_59_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_67_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_67_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_75_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_75_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_11_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_11_sg1 <= 17'b0;
      else_7_if_1_div_9cyc_st_3 <= 4'b0;
      delta_conc_2_tmp_mut_11_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_11_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_19_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_19_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_27_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_27_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_35_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_35_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_43_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_43_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_51_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_51_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_59_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_59_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_67_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_67_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_75_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_75_sg1 <= 17'b0;
      else_7_else_1_if_div_9cyc_st_3 <= 4'b0;
      delta_conc_3_tmp_mut_11_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_11_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_19_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_19_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_27_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_27_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_35_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_35_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_43_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_43_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_51_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_51_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_59_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_59_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_67_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_67_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_75_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_75_sg1 <= 17'b0;
      else_7_else_1_else_div_9cyc_st_3 <= 4'b0;
      else_7_else_1_equal_svs_st_3 <= 1'b0;
      else_7_equal_svs_st_3 <= 1'b0;
      max_sg1_lpi_dfm_3_st_3 <= 16'b0;
      if_7_equal_svs_st_3 <= 1'b0;
      max_conc_4_tmp_mut_18_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_18_sg1 <= 16'b0;
      max_conc_4_tmp_mut_26_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_26_sg1 <= 16'b0;
      max_conc_4_tmp_mut_34_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_34_sg1 <= 16'b0;
      max_conc_4_tmp_mut_42_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_42_sg1 <= 16'b0;
      max_conc_4_tmp_mut_50_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_50_sg1 <= 16'b0;
      max_conc_4_tmp_mut_58_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_58_sg1 <= 16'b0;
      max_conc_4_tmp_mut_66_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_66_sg1 <= 16'b0;
      max_conc_4_tmp_mut_74_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_74_sg1 <= 16'b0;
      max_conc_4_tmp_mut_10_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_10_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_2 <= 4'b0;
      delta_conc_1_tmp_mut_18_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_18_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_26_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_26_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_34_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_34_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_42_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_42_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_50_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_50_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_58_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_58_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_66_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_66_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_74_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_74_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_10_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_10_sg1 <= 17'b0;
      else_7_if_1_div_9cyc_st_2 <= 4'b0;
      delta_conc_2_tmp_mut_10_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_10_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_18_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_18_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_26_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_26_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_34_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_34_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_42_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_42_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_50_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_50_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_58_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_58_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_66_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_66_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_74_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_74_sg1 <= 17'b0;
      else_7_else_1_if_div_9cyc_st_2 <= 4'b0;
      delta_conc_3_tmp_mut_10_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_10_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_18_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_18_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_26_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_26_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_34_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_34_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_42_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_42_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_50_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_50_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_58_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_58_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_66_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_66_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_74_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_74_sg1 <= 17'b0;
      else_7_else_1_else_div_9cyc_st_2 <= 4'b0;
      else_7_else_1_equal_svs_st_2 <= 1'b0;
      else_7_equal_svs_st_2 <= 1'b0;
      max_sg1_lpi_dfm_3_st_2 <= 16'b0;
      if_7_equal_svs_st_2 <= 1'b0;
      max_conc_4_tmp_mut_17_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_17_sg1 <= 16'b0;
      max_conc_4_tmp_mut_25_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_25_sg1 <= 16'b0;
      max_conc_4_tmp_mut_33_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_33_sg1 <= 16'b0;
      max_conc_4_tmp_mut_41_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_41_sg1 <= 16'b0;
      max_conc_4_tmp_mut_49_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_49_sg1 <= 16'b0;
      max_conc_4_tmp_mut_57_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_57_sg1 <= 16'b0;
      max_conc_4_tmp_mut_65_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_65_sg1 <= 16'b0;
      max_conc_4_tmp_mut_73_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_73_sg1 <= 16'b0;
      max_conc_4_tmp_mut_9_sg1 <= 16'b0;
      else_7_if_conc_tmp_mut_9_sg1 <= 16'b0;
      else_7_if_div_9cyc_st_1 <= 4'b0;
      delta_conc_1_tmp_mut_17_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_17_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_25_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_25_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_33_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_33_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_41_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_41_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_49_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_49_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_57_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_57_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_65_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_65_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_73_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_73_sg1 <= 17'b0;
      delta_conc_1_tmp_mut_9_sg1 <= 16'b0;
      else_7_if_1_conc_tmp_mut_9_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_9_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_9_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_17_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_17_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_25_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_25_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_33_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_33_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_41_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_41_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_49_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_49_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_57_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_57_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_65_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_65_sg1 <= 17'b0;
      delta_conc_2_tmp_mut_73_sg1 <= 16'b0;
      else_7_else_1_if_conc_tmp_mut_73_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_9_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_9_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_17_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_17_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_25_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_25_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_33_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_33_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_41_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_41_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_49_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_49_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_57_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_57_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_65_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_65_sg1 <= 17'b0;
      delta_conc_3_tmp_mut_73_sg1 <= 16'b0;
      else_7_else_1_else_conc_tmp_mut_73_sg1 <= 17'b0;
      else_7_equal_svs_st_1 <= 1'b0;
      max_sg1_lpi_dfm_3_st_1 <= 16'b0;
      if_7_equal_svs_st_1 <= 1'b0;
      else_7_if_div_9cyc <= 4'b0;
      else_7_if_1_div_9cyc <= 4'b0;
      else_7_else_1_if_div_9cyc <= 4'b0;
      else_7_else_1_else_div_9cyc <= 4'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      main_stage_0_7 <= 1'b0;
      main_stage_0_8 <= 1'b0;
      main_stage_0_9 <= 1'b0;
      main_stage_0_10 <= 1'b0;
      else_7_if_div_9cyc_st <= 4'b0;
      slc_3_itm_8 <= 15'b0;
      else_7_and_5_itm_8 <= 1'b0;
      unequal_tmp_8 <= 1'b0;
      slc_3_itm_7 <= 15'b0;
      else_7_and_5_itm_7 <= 1'b0;
      unequal_tmp_7 <= 1'b0;
      slc_3_itm_6 <= 15'b0;
      else_7_and_5_itm_6 <= 1'b0;
      unequal_tmp_6 <= 1'b0;
      slc_3_itm_5 <= 15'b0;
      else_7_and_5_itm_5 <= 1'b0;
      unequal_tmp_5 <= 1'b0;
      slc_3_itm_4 <= 15'b0;
      else_7_and_5_itm_4 <= 1'b0;
      unequal_tmp_4 <= 1'b0;
      slc_3_itm_3 <= 15'b0;
      else_7_and_5_itm_3 <= 1'b0;
      unequal_tmp_3 <= 1'b0;
      slc_3_itm_2 <= 15'b0;
      else_7_and_5_itm_2 <= 1'b0;
      unequal_tmp_2 <= 1'b0;
      slc_3_itm_1 <= 15'b0;
      else_7_and_5_itm_1 <= 1'b0;
      unequal_tmp_1 <= 1'b0;
      else_7_else_1_equal_svs_1 <= 1'b0;
      reg_div_mgc_div_28_b_tmp <= 16'b0;
      reg_div_mgc_div_28_a_tmp <= 16'b0;
      reg_div_mgc_div_29_b_tmp <= 16'b0;
      reg_div_mgc_div_29_a_tmp <= 16'b0;
      reg_div_mgc_div_30_b_tmp <= 16'b0;
      reg_div_mgc_div_30_a_tmp <= 16'b0;
      reg_div_mgc_div_31_b_tmp <= 16'b0;
      reg_div_mgc_div_31_a_tmp <= 16'b0;
      reg_div_mgc_div_32_b_tmp <= 16'b0;
      reg_div_mgc_div_32_a_tmp <= 16'b0;
      reg_div_mgc_div_33_b_tmp <= 16'b0;
      reg_div_mgc_div_33_a_tmp <= 16'b0;
      reg_div_mgc_div_34_b_tmp <= 16'b0;
      reg_div_mgc_div_34_a_tmp <= 16'b0;
      reg_div_mgc_div_35_b_tmp <= 16'b0;
      reg_div_mgc_div_35_a_tmp <= 16'b0;
      reg_div_mgc_div_27_b_tmp <= 16'b0;
      reg_div_mgc_div_27_a_tmp <= 16'b0;
      reg_div_mgc_div_19_b_tmp <= 16'b0;
      reg_div_mgc_div_19_a_tmp <= 17'b0;
      reg_div_mgc_div_20_b_tmp <= 16'b0;
      reg_div_mgc_div_20_a_tmp <= 17'b0;
      reg_div_mgc_div_21_b_tmp <= 16'b0;
      reg_div_mgc_div_21_a_tmp <= 17'b0;
      reg_div_mgc_div_22_b_tmp <= 16'b0;
      reg_div_mgc_div_22_a_tmp <= 17'b0;
      reg_div_mgc_div_23_b_tmp <= 16'b0;
      reg_div_mgc_div_23_a_tmp <= 17'b0;
      reg_div_mgc_div_24_b_tmp <= 16'b0;
      reg_div_mgc_div_24_a_tmp <= 17'b0;
      reg_div_mgc_div_25_b_tmp <= 16'b0;
      reg_div_mgc_div_25_a_tmp <= 17'b0;
      reg_div_mgc_div_26_b_tmp <= 16'b0;
      reg_div_mgc_div_26_a_tmp <= 17'b0;
      reg_div_mgc_div_b_tmp <= 16'b0;
      reg_div_mgc_div_a_tmp <= 17'b0;
      reg_div_mgc_div_10_b_tmp <= 16'b0;
      reg_div_mgc_div_10_a_tmp <= 17'b0;
      reg_div_mgc_div_11_b_tmp <= 16'b0;
      reg_div_mgc_div_11_a_tmp <= 17'b0;
      reg_div_mgc_div_12_b_tmp <= 16'b0;
      reg_div_mgc_div_12_a_tmp <= 17'b0;
      reg_div_mgc_div_13_b_tmp <= 16'b0;
      reg_div_mgc_div_13_a_tmp <= 17'b0;
      reg_div_mgc_div_14_b_tmp <= 16'b0;
      reg_div_mgc_div_14_a_tmp <= 17'b0;
      reg_div_mgc_div_15_b_tmp <= 16'b0;
      reg_div_mgc_div_15_a_tmp <= 17'b0;
      reg_div_mgc_div_16_b_tmp <= 16'b0;
      reg_div_mgc_div_16_a_tmp <= 17'b0;
      reg_div_mgc_div_17_b_tmp <= 16'b0;
      reg_div_mgc_div_17_a_tmp <= 17'b0;
      reg_div_mgc_div_18_b_tmp <= 16'b0;
      reg_div_mgc_div_18_a_tmp <= 17'b0;
      reg_div_mgc_div_1_b_tmp <= 16'b0;
      reg_div_mgc_div_1_a_tmp <= 17'b0;
      reg_div_mgc_div_2_b_tmp <= 16'b0;
      reg_div_mgc_div_2_a_tmp <= 17'b0;
      reg_div_mgc_div_3_b_tmp <= 16'b0;
      reg_div_mgc_div_3_a_tmp <= 17'b0;
      reg_div_mgc_div_4_b_tmp <= 16'b0;
      reg_div_mgc_div_4_a_tmp <= 17'b0;
      reg_div_mgc_div_5_b_tmp <= 16'b0;
      reg_div_mgc_div_5_a_tmp <= 17'b0;
      reg_div_mgc_div_6_b_tmp <= 16'b0;
      reg_div_mgc_div_6_a_tmp <= 17'b0;
      reg_div_mgc_div_7_b_tmp <= 16'b0;
      reg_div_mgc_div_7_a_tmp <= 17'b0;
      reg_div_mgc_div_8_b_tmp <= 16'b0;
      reg_div_mgc_div_8_a_tmp <= 17'b0;
      reg_div_mgc_div_9_b_tmp <= 16'b0;
      reg_div_mgc_div_9_a_tmp <= 17'b0;
    end
    else begin
      V_OUT_rsc_mgc_out_stdreg_d <= MUX_v_32_2_2({V_OUT_rsc_mgc_out_stdreg_d , ({{17{slc_3_itm_9[14]}},
          slc_3_itm_9})}, main_stage_0_10);
      S_OUT_rsc_mgc_out_stdreg_d <= MUX_v_32_2_2({S_OUT_rsc_mgc_out_stdreg_d , ({(signext_30_21(conv_s2u_42_21(conv_s2s_16_21((MUX1HOT_v_16_10_2({(div_mgc_div_28_z[31:16])
          , (div_mgc_div_29_z[31:16]) , (div_mgc_div_30_z[31:16]) , (div_mgc_div_31_z[31:16])
          , (div_mgc_div_32_z[31:16]) , (div_mgc_div_33_z[31:16]) , (div_mgc_div_34_z[31:16])
          , (div_mgc_div_35_z[31:16]) , (div_mgc_div_27_z[31:16]) , else_7_if_div_tmp_duc_sg1},
          {(or_303_cse & and_dcpl_2742 & and_dcpl_2741) , (or_303_cse & and_dcpl_2746
          & and_dcpl_2741) , (or_303_cse & and_dcpl_2742 & and_dcpl_2749) , (or_303_cse
          & and_dcpl_2746 & and_dcpl_2749) , (or_303_cse & and_dcpl_2742 & and_dcpl_2757)
          , (or_303_cse & and_dcpl_2746 & and_dcpl_2757) , (or_303_cse & and_dcpl_2742
          & and_dcpl_2765) , (or_303_cse & and_dcpl_2746 & and_dcpl_2765) , (or_303_cse
          & (else_7_if_div_9cyc_st_9[3]) & (~ (else_7_if_div_9cyc_st_9[0])) & and_dcpl_2741)
          , or_tmp_4})) & ({{15{unequal_tmp_9}}, unequal_tmp_9}) & (signext_16_1(~
          if_7_equal_svs_9))) * 21'b11001))) , 2'b0})}, main_stage_0_10);
      H_OUT_rsc_mgc_out_stdreg_d <= MUX_v_32_2_2({H_OUT_rsc_mgc_out_stdreg_d , (signext_32_16({((MUX_v_13_2_2({(else_7_acc_2_psp_sg1_sva_1[15:3])
          , (({1'b1 , (else_7_acc_2_itm[28:17])}) + 13'b101101)}, else_7_acc_2_psp_sg1_sva_1[15]))
          & (signext_13_1(~ if_7_equal_svs_9))) , ((else_7_acc_2_psp_sg1_sva_1[2:0])
          & (signext_3_1(~ if_7_equal_svs_9)))}))}, main_stage_0_10);
      else_7_acc_2_psp_sg1_sva <= MUX_v_16_2_2({else_7_acc_2_psp_sg1_sva , (else_7_acc_2_itm[29:14])},
          and_9092_cse);
      else_7_if_div_tmp_duc_sg1 <= MUX1HOT_v_16_10_2({(div_mgc_div_28_z[31:16]) ,
          (div_mgc_div_29_z[31:16]) , (div_mgc_div_30_z[31:16]) , (div_mgc_div_31_z[31:16])
          , (div_mgc_div_32_z[31:16]) , (div_mgc_div_33_z[31:16]) , (div_mgc_div_34_z[31:16])
          , (div_mgc_div_35_z[31:16]) , (div_mgc_div_27_z[31:16]) , else_7_if_div_tmp_duc_sg1},
          {(or_303_cse & and_dcpl_2780 & and_dcpl_2778) , (or_303_cse & and_dcpl_2780
          & and_dcpl_2783 & (~ (else_7_if_div_9cyc_st_9[2]))) , (or_303_cse & and_dcpl_2780
          & and_dcpl_2789 & (~ (else_7_if_div_9cyc_st_9[2]))) , (or_303_cse & and_dcpl_2780
          & and_dcpl_2795 & (~ (else_7_if_div_9cyc_st_9[2]))) , (or_303_cse & and_dcpl_2780
          & and_dcpl_2777 & (else_7_if_div_9cyc_st_9[2])) , (or_303_cse & and_dcpl_2780
          & and_dcpl_2783 & (else_7_if_div_9cyc_st_9[2])) , (or_303_cse & and_dcpl_2780
          & and_dcpl_2789 & (else_7_if_div_9cyc_st_9[2])) , (or_303_cse & and_dcpl_2780
          & and_dcpl_2795 & (else_7_if_div_9cyc_st_9[2])) , (or_303_cse & and_9092_cse
          & (else_7_if_div_9cyc_st_9[3]) & and_dcpl_2778) , (or_tmp_4 | or_dcpl_555)});
      else_7_if_div_9cyc_st_9 <= else_7_if_div_9cyc_st_8;
      h_2_sva_duc <= MUX1HOT_v_30_10_2({(div_mgc_div_19_z[29:0]) , (div_mgc_div_20_z[29:0])
          , (div_mgc_div_21_z[29:0]) , (div_mgc_div_22_z[29:0]) , (div_mgc_div_23_z[29:0])
          , (div_mgc_div_24_z[29:0]) , (div_mgc_div_25_z[29:0]) , (div_mgc_div_26_z[29:0])
          , (div_mgc_div_z[29:0]) , h_2_sva_duc}, {(and_dcpl_2863 & and_dcpl_2860)
          , (and_dcpl_2863 & and_dcpl_2865 & (~ (else_7_if_1_div_9cyc_st_9[2])))
          , (and_dcpl_2863 & and_dcpl_2871 & (~ (else_7_if_1_div_9cyc_st_9[2])))
          , (and_dcpl_2863 & and_dcpl_2877 & (~ (else_7_if_1_div_9cyc_st_9[2])))
          , (and_dcpl_2863 & and_dcpl_2859 & (else_7_if_1_div_9cyc_st_9[2])) , (and_dcpl_2863
          & and_dcpl_2865 & (else_7_if_1_div_9cyc_st_9[2])) , (and_dcpl_2863 & and_dcpl_2871
          & (else_7_if_1_div_9cyc_st_9[2])) , (and_dcpl_2863 & and_dcpl_2877 & (else_7_if_1_div_9cyc_st_9[2]))
          , (and_9092_cse & else_7_equal_svs_9 & (else_7_if_1_div_9cyc_st_9[3]) &
          and_dcpl_2860) , (and_2924_cse | or_dcpl_555 | (~ else_7_equal_svs_9))});
      else_7_if_1_div_9cyc_st_9 <= else_7_if_1_div_9cyc_st_8;
      div_sdt_2_sva_duc <= MUX1HOT_v_30_10_2({(div_mgc_div_10_z[29:0]) , (div_mgc_div_11_z[29:0])
          , (div_mgc_div_12_z[29:0]) , (div_mgc_div_13_z[29:0]) , (div_mgc_div_14_z[29:0])
          , (div_mgc_div_15_z[29:0]) , (div_mgc_div_16_z[29:0]) , (div_mgc_div_17_z[29:0])
          , (div_mgc_div_18_z[29:0]) , div_sdt_2_sva_duc}, {(and_dcpl_2993 & and_2973_cse)
          , (and_dcpl_2993 & and_2976_cse) , (and_dcpl_2993 & and_2979_cse) , (and_dcpl_2993
          & and_2982_cse) , (and_dcpl_2993 & and_2985_cse) , (and_dcpl_2993 & and_2988_cse)
          , (and_dcpl_2993 & and_2991_cse) , (and_dcpl_2993 & and_2994_cse) , (and_dcpl_2993
          & and_2997_cse) , (and_3062_cse | or_dcpl_555 | or_dcpl_564)});
      div_sdt_3_sva_duc <= MUX1HOT_v_30_10_2({(div_mgc_div_1_z[29:0]) , (div_mgc_div_2_z[29:0])
          , (div_mgc_div_3_z[29:0]) , (div_mgc_div_4_z[29:0]) , (div_mgc_div_5_z[29:0])
          , (div_mgc_div_6_z[29:0]) , (div_mgc_div_7_z[29:0]) , (div_mgc_div_8_z[29:0])
          , (div_mgc_div_9_z[29:0]) , div_sdt_3_sva_duc}, {(and_dcpl_3085 & and_3065_cse)
          , (and_dcpl_3085 & and_3068_cse) , (and_dcpl_3085 & and_3071_cse) , (and_dcpl_3085
          & and_3074_cse) , (and_dcpl_3085 & and_3077_cse) , (and_dcpl_3085 & and_3080_cse)
          , (and_dcpl_3085 & and_3083_cse) , (and_dcpl_3085 & and_3086_cse) , (and_dcpl_3085
          & and_3089_cse) , (and_3154_cse | or_dcpl_555 | else_7_equal_svs_9 | else_7_else_1_equal_svs_st_9)});
      else_7_else_1_if_div_9cyc_st_9 <= else_7_else_1_if_div_9cyc_st_8;
      else_7_else_1_else_div_9cyc_st_9 <= else_7_else_1_else_div_9cyc_st_8;
      else_7_else_1_equal_svs_st_9 <= else_7_else_1_equal_svs_st_8;
      else_7_and_5_itm_9 <= else_7_and_5_itm_8;
      else_7_equal_svs_9 <= else_7_equal_svs_st_8;
      unequal_tmp_9 <= unequal_tmp_8;
      max_sg1_lpi_dfm_3_st_9 <= max_sg1_lpi_dfm_3_st_8;
      slc_3_itm_9 <= slc_3_itm_8;
      if_7_equal_svs_9 <= if_7_equal_svs_st_8;
      max_conc_4_tmp_mut_24_sg1 <= max_conc_4_tmp_mut_23_sg1;
      else_7_if_conc_tmp_mut_24_sg1 <= else_7_if_conc_tmp_mut_23_sg1;
      max_conc_4_tmp_mut_32_sg1 <= max_conc_4_tmp_mut_31_sg1;
      else_7_if_conc_tmp_mut_32_sg1 <= else_7_if_conc_tmp_mut_31_sg1;
      max_conc_4_tmp_mut_40_sg1 <= max_conc_4_tmp_mut_39_sg1;
      else_7_if_conc_tmp_mut_40_sg1 <= else_7_if_conc_tmp_mut_39_sg1;
      max_conc_4_tmp_mut_48_sg1 <= max_conc_4_tmp_mut_47_sg1;
      else_7_if_conc_tmp_mut_48_sg1 <= else_7_if_conc_tmp_mut_47_sg1;
      max_conc_4_tmp_mut_56_sg1 <= max_conc_4_tmp_mut_55_sg1;
      else_7_if_conc_tmp_mut_56_sg1 <= else_7_if_conc_tmp_mut_55_sg1;
      max_conc_4_tmp_mut_64_sg1 <= max_conc_4_tmp_mut_63_sg1;
      else_7_if_conc_tmp_mut_64_sg1 <= else_7_if_conc_tmp_mut_63_sg1;
      max_conc_4_tmp_mut_72_sg1 <= max_conc_4_tmp_mut_71_sg1;
      else_7_if_conc_tmp_mut_72_sg1 <= else_7_if_conc_tmp_mut_71_sg1;
      max_conc_4_tmp_mut_80_sg1 <= max_conc_4_tmp_mut_79_sg1;
      else_7_if_conc_tmp_mut_80_sg1 <= else_7_if_conc_tmp_mut_79_sg1;
      max_conc_4_tmp_mut_16_sg1 <= max_conc_4_tmp_mut_15_sg1;
      else_7_if_conc_tmp_mut_16_sg1 <= else_7_if_conc_tmp_mut_15_sg1;
      else_7_if_div_9cyc_st_8 <= else_7_if_div_9cyc_st_7;
      delta_conc_1_tmp_mut_24_sg1 <= delta_conc_1_tmp_mut_23_sg1;
      else_7_if_1_conc_tmp_mut_24_sg1 <= else_7_if_1_conc_tmp_mut_23_sg1;
      delta_conc_1_tmp_mut_32_sg1 <= delta_conc_1_tmp_mut_31_sg1;
      else_7_if_1_conc_tmp_mut_32_sg1 <= else_7_if_1_conc_tmp_mut_31_sg1;
      delta_conc_1_tmp_mut_40_sg1 <= delta_conc_1_tmp_mut_39_sg1;
      else_7_if_1_conc_tmp_mut_40_sg1 <= else_7_if_1_conc_tmp_mut_39_sg1;
      delta_conc_1_tmp_mut_48_sg1 <= delta_conc_1_tmp_mut_47_sg1;
      else_7_if_1_conc_tmp_mut_48_sg1 <= else_7_if_1_conc_tmp_mut_47_sg1;
      delta_conc_1_tmp_mut_56_sg1 <= delta_conc_1_tmp_mut_55_sg1;
      else_7_if_1_conc_tmp_mut_56_sg1 <= else_7_if_1_conc_tmp_mut_55_sg1;
      delta_conc_1_tmp_mut_64_sg1 <= delta_conc_1_tmp_mut_63_sg1;
      else_7_if_1_conc_tmp_mut_64_sg1 <= else_7_if_1_conc_tmp_mut_63_sg1;
      delta_conc_1_tmp_mut_72_sg1 <= delta_conc_1_tmp_mut_71_sg1;
      else_7_if_1_conc_tmp_mut_72_sg1 <= else_7_if_1_conc_tmp_mut_71_sg1;
      delta_conc_1_tmp_mut_80_sg1 <= delta_conc_1_tmp_mut_79_sg1;
      else_7_if_1_conc_tmp_mut_80_sg1 <= else_7_if_1_conc_tmp_mut_79_sg1;
      delta_conc_1_tmp_mut_16_sg1 <= delta_conc_1_tmp_mut_15_sg1;
      else_7_if_1_conc_tmp_mut_16_sg1 <= else_7_if_1_conc_tmp_mut_15_sg1;
      else_7_if_1_div_9cyc_st_8 <= else_7_if_1_div_9cyc_st_7;
      delta_conc_2_tmp_mut_16_sg1 <= delta_conc_2_tmp_mut_15_sg1;
      else_7_else_1_if_conc_tmp_mut_16_sg1 <= else_7_else_1_if_conc_tmp_mut_15_sg1;
      delta_conc_2_tmp_mut_24_sg1 <= delta_conc_2_tmp_mut_23_sg1;
      else_7_else_1_if_conc_tmp_mut_24_sg1 <= else_7_else_1_if_conc_tmp_mut_23_sg1;
      delta_conc_2_tmp_mut_32_sg1 <= delta_conc_2_tmp_mut_31_sg1;
      else_7_else_1_if_conc_tmp_mut_32_sg1 <= else_7_else_1_if_conc_tmp_mut_31_sg1;
      delta_conc_2_tmp_mut_40_sg1 <= delta_conc_2_tmp_mut_39_sg1;
      else_7_else_1_if_conc_tmp_mut_40_sg1 <= else_7_else_1_if_conc_tmp_mut_39_sg1;
      delta_conc_2_tmp_mut_48_sg1 <= delta_conc_2_tmp_mut_47_sg1;
      else_7_else_1_if_conc_tmp_mut_48_sg1 <= else_7_else_1_if_conc_tmp_mut_47_sg1;
      delta_conc_2_tmp_mut_56_sg1 <= delta_conc_2_tmp_mut_55_sg1;
      else_7_else_1_if_conc_tmp_mut_56_sg1 <= else_7_else_1_if_conc_tmp_mut_55_sg1;
      delta_conc_2_tmp_mut_64_sg1 <= delta_conc_2_tmp_mut_63_sg1;
      else_7_else_1_if_conc_tmp_mut_64_sg1 <= else_7_else_1_if_conc_tmp_mut_63_sg1;
      delta_conc_2_tmp_mut_72_sg1 <= delta_conc_2_tmp_mut_71_sg1;
      else_7_else_1_if_conc_tmp_mut_72_sg1 <= else_7_else_1_if_conc_tmp_mut_71_sg1;
      delta_conc_2_tmp_mut_80_sg1 <= delta_conc_2_tmp_mut_79_sg1;
      else_7_else_1_if_conc_tmp_mut_80_sg1 <= else_7_else_1_if_conc_tmp_mut_79_sg1;
      else_7_else_1_if_div_9cyc_st_8 <= else_7_else_1_if_div_9cyc_st_7;
      delta_conc_3_tmp_mut_16_sg1 <= delta_conc_3_tmp_mut_15_sg1;
      else_7_else_1_else_conc_tmp_mut_16_sg1 <= else_7_else_1_else_conc_tmp_mut_15_sg1;
      delta_conc_3_tmp_mut_24_sg1 <= delta_conc_3_tmp_mut_23_sg1;
      else_7_else_1_else_conc_tmp_mut_24_sg1 <= else_7_else_1_else_conc_tmp_mut_23_sg1;
      delta_conc_3_tmp_mut_32_sg1 <= delta_conc_3_tmp_mut_31_sg1;
      else_7_else_1_else_conc_tmp_mut_32_sg1 <= else_7_else_1_else_conc_tmp_mut_31_sg1;
      delta_conc_3_tmp_mut_40_sg1 <= delta_conc_3_tmp_mut_39_sg1;
      else_7_else_1_else_conc_tmp_mut_40_sg1 <= else_7_else_1_else_conc_tmp_mut_39_sg1;
      delta_conc_3_tmp_mut_48_sg1 <= delta_conc_3_tmp_mut_47_sg1;
      else_7_else_1_else_conc_tmp_mut_48_sg1 <= else_7_else_1_else_conc_tmp_mut_47_sg1;
      delta_conc_3_tmp_mut_56_sg1 <= delta_conc_3_tmp_mut_55_sg1;
      else_7_else_1_else_conc_tmp_mut_56_sg1 <= else_7_else_1_else_conc_tmp_mut_55_sg1;
      delta_conc_3_tmp_mut_64_sg1 <= delta_conc_3_tmp_mut_63_sg1;
      else_7_else_1_else_conc_tmp_mut_64_sg1 <= else_7_else_1_else_conc_tmp_mut_63_sg1;
      delta_conc_3_tmp_mut_72_sg1 <= delta_conc_3_tmp_mut_71_sg1;
      else_7_else_1_else_conc_tmp_mut_72_sg1 <= else_7_else_1_else_conc_tmp_mut_71_sg1;
      delta_conc_3_tmp_mut_80_sg1 <= delta_conc_3_tmp_mut_79_sg1;
      else_7_else_1_else_conc_tmp_mut_80_sg1 <= else_7_else_1_else_conc_tmp_mut_79_sg1;
      else_7_else_1_else_div_9cyc_st_8 <= else_7_else_1_else_div_9cyc_st_7;
      else_7_else_1_equal_svs_st_8 <= else_7_else_1_equal_svs_st_7;
      else_7_equal_svs_st_8 <= else_7_equal_svs_st_7;
      max_sg1_lpi_dfm_3_st_8 <= max_sg1_lpi_dfm_3_st_7;
      if_7_equal_svs_st_8 <= if_7_equal_svs_st_7;
      max_conc_4_tmp_mut_23_sg1 <= max_conc_4_tmp_mut_22_sg1;
      else_7_if_conc_tmp_mut_23_sg1 <= else_7_if_conc_tmp_mut_22_sg1;
      max_conc_4_tmp_mut_31_sg1 <= max_conc_4_tmp_mut_30_sg1;
      else_7_if_conc_tmp_mut_31_sg1 <= else_7_if_conc_tmp_mut_30_sg1;
      max_conc_4_tmp_mut_39_sg1 <= max_conc_4_tmp_mut_38_sg1;
      else_7_if_conc_tmp_mut_39_sg1 <= else_7_if_conc_tmp_mut_38_sg1;
      max_conc_4_tmp_mut_47_sg1 <= max_conc_4_tmp_mut_46_sg1;
      else_7_if_conc_tmp_mut_47_sg1 <= else_7_if_conc_tmp_mut_46_sg1;
      max_conc_4_tmp_mut_55_sg1 <= max_conc_4_tmp_mut_54_sg1;
      else_7_if_conc_tmp_mut_55_sg1 <= else_7_if_conc_tmp_mut_54_sg1;
      max_conc_4_tmp_mut_63_sg1 <= max_conc_4_tmp_mut_62_sg1;
      else_7_if_conc_tmp_mut_63_sg1 <= else_7_if_conc_tmp_mut_62_sg1;
      max_conc_4_tmp_mut_71_sg1 <= max_conc_4_tmp_mut_70_sg1;
      else_7_if_conc_tmp_mut_71_sg1 <= else_7_if_conc_tmp_mut_70_sg1;
      max_conc_4_tmp_mut_79_sg1 <= max_conc_4_tmp_mut_78_sg1;
      else_7_if_conc_tmp_mut_79_sg1 <= else_7_if_conc_tmp_mut_78_sg1;
      max_conc_4_tmp_mut_15_sg1 <= max_conc_4_tmp_mut_14_sg1;
      else_7_if_conc_tmp_mut_15_sg1 <= else_7_if_conc_tmp_mut_14_sg1;
      else_7_if_div_9cyc_st_7 <= else_7_if_div_9cyc_st_6;
      delta_conc_1_tmp_mut_23_sg1 <= delta_conc_1_tmp_mut_22_sg1;
      else_7_if_1_conc_tmp_mut_23_sg1 <= else_7_if_1_conc_tmp_mut_22_sg1;
      delta_conc_1_tmp_mut_31_sg1 <= delta_conc_1_tmp_mut_30_sg1;
      else_7_if_1_conc_tmp_mut_31_sg1 <= else_7_if_1_conc_tmp_mut_30_sg1;
      delta_conc_1_tmp_mut_39_sg1 <= delta_conc_1_tmp_mut_38_sg1;
      else_7_if_1_conc_tmp_mut_39_sg1 <= else_7_if_1_conc_tmp_mut_38_sg1;
      delta_conc_1_tmp_mut_47_sg1 <= delta_conc_1_tmp_mut_46_sg1;
      else_7_if_1_conc_tmp_mut_47_sg1 <= else_7_if_1_conc_tmp_mut_46_sg1;
      delta_conc_1_tmp_mut_55_sg1 <= delta_conc_1_tmp_mut_54_sg1;
      else_7_if_1_conc_tmp_mut_55_sg1 <= else_7_if_1_conc_tmp_mut_54_sg1;
      delta_conc_1_tmp_mut_63_sg1 <= delta_conc_1_tmp_mut_62_sg1;
      else_7_if_1_conc_tmp_mut_63_sg1 <= else_7_if_1_conc_tmp_mut_62_sg1;
      delta_conc_1_tmp_mut_71_sg1 <= delta_conc_1_tmp_mut_70_sg1;
      else_7_if_1_conc_tmp_mut_71_sg1 <= else_7_if_1_conc_tmp_mut_70_sg1;
      delta_conc_1_tmp_mut_79_sg1 <= delta_conc_1_tmp_mut_78_sg1;
      else_7_if_1_conc_tmp_mut_79_sg1 <= else_7_if_1_conc_tmp_mut_78_sg1;
      delta_conc_1_tmp_mut_15_sg1 <= delta_conc_1_tmp_mut_14_sg1;
      else_7_if_1_conc_tmp_mut_15_sg1 <= else_7_if_1_conc_tmp_mut_14_sg1;
      else_7_if_1_div_9cyc_st_7 <= else_7_if_1_div_9cyc_st_6;
      delta_conc_2_tmp_mut_15_sg1 <= delta_conc_2_tmp_mut_14_sg1;
      else_7_else_1_if_conc_tmp_mut_15_sg1 <= else_7_else_1_if_conc_tmp_mut_14_sg1;
      delta_conc_2_tmp_mut_23_sg1 <= delta_conc_2_tmp_mut_22_sg1;
      else_7_else_1_if_conc_tmp_mut_23_sg1 <= else_7_else_1_if_conc_tmp_mut_22_sg1;
      delta_conc_2_tmp_mut_31_sg1 <= delta_conc_2_tmp_mut_30_sg1;
      else_7_else_1_if_conc_tmp_mut_31_sg1 <= else_7_else_1_if_conc_tmp_mut_30_sg1;
      delta_conc_2_tmp_mut_39_sg1 <= delta_conc_2_tmp_mut_38_sg1;
      else_7_else_1_if_conc_tmp_mut_39_sg1 <= else_7_else_1_if_conc_tmp_mut_38_sg1;
      delta_conc_2_tmp_mut_47_sg1 <= delta_conc_2_tmp_mut_46_sg1;
      else_7_else_1_if_conc_tmp_mut_47_sg1 <= else_7_else_1_if_conc_tmp_mut_46_sg1;
      delta_conc_2_tmp_mut_55_sg1 <= delta_conc_2_tmp_mut_54_sg1;
      else_7_else_1_if_conc_tmp_mut_55_sg1 <= else_7_else_1_if_conc_tmp_mut_54_sg1;
      delta_conc_2_tmp_mut_63_sg1 <= delta_conc_2_tmp_mut_62_sg1;
      else_7_else_1_if_conc_tmp_mut_63_sg1 <= else_7_else_1_if_conc_tmp_mut_62_sg1;
      delta_conc_2_tmp_mut_71_sg1 <= delta_conc_2_tmp_mut_70_sg1;
      else_7_else_1_if_conc_tmp_mut_71_sg1 <= else_7_else_1_if_conc_tmp_mut_70_sg1;
      delta_conc_2_tmp_mut_79_sg1 <= delta_conc_2_tmp_mut_78_sg1;
      else_7_else_1_if_conc_tmp_mut_79_sg1 <= else_7_else_1_if_conc_tmp_mut_78_sg1;
      else_7_else_1_if_div_9cyc_st_7 <= else_7_else_1_if_div_9cyc_st_6;
      delta_conc_3_tmp_mut_15_sg1 <= delta_conc_3_tmp_mut_14_sg1;
      else_7_else_1_else_conc_tmp_mut_15_sg1 <= else_7_else_1_else_conc_tmp_mut_14_sg1;
      delta_conc_3_tmp_mut_23_sg1 <= delta_conc_3_tmp_mut_22_sg1;
      else_7_else_1_else_conc_tmp_mut_23_sg1 <= else_7_else_1_else_conc_tmp_mut_22_sg1;
      delta_conc_3_tmp_mut_31_sg1 <= delta_conc_3_tmp_mut_30_sg1;
      else_7_else_1_else_conc_tmp_mut_31_sg1 <= else_7_else_1_else_conc_tmp_mut_30_sg1;
      delta_conc_3_tmp_mut_39_sg1 <= delta_conc_3_tmp_mut_38_sg1;
      else_7_else_1_else_conc_tmp_mut_39_sg1 <= else_7_else_1_else_conc_tmp_mut_38_sg1;
      delta_conc_3_tmp_mut_47_sg1 <= delta_conc_3_tmp_mut_46_sg1;
      else_7_else_1_else_conc_tmp_mut_47_sg1 <= else_7_else_1_else_conc_tmp_mut_46_sg1;
      delta_conc_3_tmp_mut_55_sg1 <= delta_conc_3_tmp_mut_54_sg1;
      else_7_else_1_else_conc_tmp_mut_55_sg1 <= else_7_else_1_else_conc_tmp_mut_54_sg1;
      delta_conc_3_tmp_mut_63_sg1 <= delta_conc_3_tmp_mut_62_sg1;
      else_7_else_1_else_conc_tmp_mut_63_sg1 <= else_7_else_1_else_conc_tmp_mut_62_sg1;
      delta_conc_3_tmp_mut_71_sg1 <= delta_conc_3_tmp_mut_70_sg1;
      else_7_else_1_else_conc_tmp_mut_71_sg1 <= else_7_else_1_else_conc_tmp_mut_70_sg1;
      delta_conc_3_tmp_mut_79_sg1 <= delta_conc_3_tmp_mut_78_sg1;
      else_7_else_1_else_conc_tmp_mut_79_sg1 <= else_7_else_1_else_conc_tmp_mut_78_sg1;
      else_7_else_1_else_div_9cyc_st_7 <= else_7_else_1_else_div_9cyc_st_6;
      else_7_else_1_equal_svs_st_7 <= else_7_else_1_equal_svs_st_6;
      else_7_equal_svs_st_7 <= else_7_equal_svs_st_6;
      max_sg1_lpi_dfm_3_st_7 <= max_sg1_lpi_dfm_3_st_6;
      if_7_equal_svs_st_7 <= if_7_equal_svs_st_6;
      max_conc_4_tmp_mut_22_sg1 <= max_conc_4_tmp_mut_21_sg1;
      else_7_if_conc_tmp_mut_22_sg1 <= else_7_if_conc_tmp_mut_21_sg1;
      max_conc_4_tmp_mut_30_sg1 <= max_conc_4_tmp_mut_29_sg1;
      else_7_if_conc_tmp_mut_30_sg1 <= else_7_if_conc_tmp_mut_29_sg1;
      max_conc_4_tmp_mut_38_sg1 <= max_conc_4_tmp_mut_37_sg1;
      else_7_if_conc_tmp_mut_38_sg1 <= else_7_if_conc_tmp_mut_37_sg1;
      max_conc_4_tmp_mut_46_sg1 <= max_conc_4_tmp_mut_45_sg1;
      else_7_if_conc_tmp_mut_46_sg1 <= else_7_if_conc_tmp_mut_45_sg1;
      max_conc_4_tmp_mut_54_sg1 <= max_conc_4_tmp_mut_53_sg1;
      else_7_if_conc_tmp_mut_54_sg1 <= else_7_if_conc_tmp_mut_53_sg1;
      max_conc_4_tmp_mut_62_sg1 <= max_conc_4_tmp_mut_61_sg1;
      else_7_if_conc_tmp_mut_62_sg1 <= else_7_if_conc_tmp_mut_61_sg1;
      max_conc_4_tmp_mut_70_sg1 <= max_conc_4_tmp_mut_69_sg1;
      else_7_if_conc_tmp_mut_70_sg1 <= else_7_if_conc_tmp_mut_69_sg1;
      max_conc_4_tmp_mut_78_sg1 <= max_conc_4_tmp_mut_77_sg1;
      else_7_if_conc_tmp_mut_78_sg1 <= else_7_if_conc_tmp_mut_77_sg1;
      max_conc_4_tmp_mut_14_sg1 <= max_conc_4_tmp_mut_13_sg1;
      else_7_if_conc_tmp_mut_14_sg1 <= else_7_if_conc_tmp_mut_13_sg1;
      else_7_if_div_9cyc_st_6 <= else_7_if_div_9cyc_st_5;
      delta_conc_1_tmp_mut_22_sg1 <= delta_conc_1_tmp_mut_21_sg1;
      else_7_if_1_conc_tmp_mut_22_sg1 <= else_7_if_1_conc_tmp_mut_21_sg1;
      delta_conc_1_tmp_mut_30_sg1 <= delta_conc_1_tmp_mut_29_sg1;
      else_7_if_1_conc_tmp_mut_30_sg1 <= else_7_if_1_conc_tmp_mut_29_sg1;
      delta_conc_1_tmp_mut_38_sg1 <= delta_conc_1_tmp_mut_37_sg1;
      else_7_if_1_conc_tmp_mut_38_sg1 <= else_7_if_1_conc_tmp_mut_37_sg1;
      delta_conc_1_tmp_mut_46_sg1 <= delta_conc_1_tmp_mut_45_sg1;
      else_7_if_1_conc_tmp_mut_46_sg1 <= else_7_if_1_conc_tmp_mut_45_sg1;
      delta_conc_1_tmp_mut_54_sg1 <= delta_conc_1_tmp_mut_53_sg1;
      else_7_if_1_conc_tmp_mut_54_sg1 <= else_7_if_1_conc_tmp_mut_53_sg1;
      delta_conc_1_tmp_mut_62_sg1 <= delta_conc_1_tmp_mut_61_sg1;
      else_7_if_1_conc_tmp_mut_62_sg1 <= else_7_if_1_conc_tmp_mut_61_sg1;
      delta_conc_1_tmp_mut_70_sg1 <= delta_conc_1_tmp_mut_69_sg1;
      else_7_if_1_conc_tmp_mut_70_sg1 <= else_7_if_1_conc_tmp_mut_69_sg1;
      delta_conc_1_tmp_mut_78_sg1 <= delta_conc_1_tmp_mut_77_sg1;
      else_7_if_1_conc_tmp_mut_78_sg1 <= else_7_if_1_conc_tmp_mut_77_sg1;
      delta_conc_1_tmp_mut_14_sg1 <= delta_conc_1_tmp_mut_13_sg1;
      else_7_if_1_conc_tmp_mut_14_sg1 <= else_7_if_1_conc_tmp_mut_13_sg1;
      else_7_if_1_div_9cyc_st_6 <= else_7_if_1_div_9cyc_st_5;
      delta_conc_2_tmp_mut_14_sg1 <= delta_conc_2_tmp_mut_13_sg1;
      else_7_else_1_if_conc_tmp_mut_14_sg1 <= else_7_else_1_if_conc_tmp_mut_13_sg1;
      delta_conc_2_tmp_mut_22_sg1 <= delta_conc_2_tmp_mut_21_sg1;
      else_7_else_1_if_conc_tmp_mut_22_sg1 <= else_7_else_1_if_conc_tmp_mut_21_sg1;
      delta_conc_2_tmp_mut_30_sg1 <= delta_conc_2_tmp_mut_29_sg1;
      else_7_else_1_if_conc_tmp_mut_30_sg1 <= else_7_else_1_if_conc_tmp_mut_29_sg1;
      delta_conc_2_tmp_mut_38_sg1 <= delta_conc_2_tmp_mut_37_sg1;
      else_7_else_1_if_conc_tmp_mut_38_sg1 <= else_7_else_1_if_conc_tmp_mut_37_sg1;
      delta_conc_2_tmp_mut_46_sg1 <= delta_conc_2_tmp_mut_45_sg1;
      else_7_else_1_if_conc_tmp_mut_46_sg1 <= else_7_else_1_if_conc_tmp_mut_45_sg1;
      delta_conc_2_tmp_mut_54_sg1 <= delta_conc_2_tmp_mut_53_sg1;
      else_7_else_1_if_conc_tmp_mut_54_sg1 <= else_7_else_1_if_conc_tmp_mut_53_sg1;
      delta_conc_2_tmp_mut_62_sg1 <= delta_conc_2_tmp_mut_61_sg1;
      else_7_else_1_if_conc_tmp_mut_62_sg1 <= else_7_else_1_if_conc_tmp_mut_61_sg1;
      delta_conc_2_tmp_mut_70_sg1 <= delta_conc_2_tmp_mut_69_sg1;
      else_7_else_1_if_conc_tmp_mut_70_sg1 <= else_7_else_1_if_conc_tmp_mut_69_sg1;
      delta_conc_2_tmp_mut_78_sg1 <= delta_conc_2_tmp_mut_77_sg1;
      else_7_else_1_if_conc_tmp_mut_78_sg1 <= else_7_else_1_if_conc_tmp_mut_77_sg1;
      else_7_else_1_if_div_9cyc_st_6 <= else_7_else_1_if_div_9cyc_st_5;
      delta_conc_3_tmp_mut_14_sg1 <= delta_conc_3_tmp_mut_13_sg1;
      else_7_else_1_else_conc_tmp_mut_14_sg1 <= else_7_else_1_else_conc_tmp_mut_13_sg1;
      delta_conc_3_tmp_mut_22_sg1 <= delta_conc_3_tmp_mut_21_sg1;
      else_7_else_1_else_conc_tmp_mut_22_sg1 <= else_7_else_1_else_conc_tmp_mut_21_sg1;
      delta_conc_3_tmp_mut_30_sg1 <= delta_conc_3_tmp_mut_29_sg1;
      else_7_else_1_else_conc_tmp_mut_30_sg1 <= else_7_else_1_else_conc_tmp_mut_29_sg1;
      delta_conc_3_tmp_mut_38_sg1 <= delta_conc_3_tmp_mut_37_sg1;
      else_7_else_1_else_conc_tmp_mut_38_sg1 <= else_7_else_1_else_conc_tmp_mut_37_sg1;
      delta_conc_3_tmp_mut_46_sg1 <= delta_conc_3_tmp_mut_45_sg1;
      else_7_else_1_else_conc_tmp_mut_46_sg1 <= else_7_else_1_else_conc_tmp_mut_45_sg1;
      delta_conc_3_tmp_mut_54_sg1 <= delta_conc_3_tmp_mut_53_sg1;
      else_7_else_1_else_conc_tmp_mut_54_sg1 <= else_7_else_1_else_conc_tmp_mut_53_sg1;
      delta_conc_3_tmp_mut_62_sg1 <= delta_conc_3_tmp_mut_61_sg1;
      else_7_else_1_else_conc_tmp_mut_62_sg1 <= else_7_else_1_else_conc_tmp_mut_61_sg1;
      delta_conc_3_tmp_mut_70_sg1 <= delta_conc_3_tmp_mut_69_sg1;
      else_7_else_1_else_conc_tmp_mut_70_sg1 <= else_7_else_1_else_conc_tmp_mut_69_sg1;
      delta_conc_3_tmp_mut_78_sg1 <= delta_conc_3_tmp_mut_77_sg1;
      else_7_else_1_else_conc_tmp_mut_78_sg1 <= else_7_else_1_else_conc_tmp_mut_77_sg1;
      else_7_else_1_else_div_9cyc_st_6 <= else_7_else_1_else_div_9cyc_st_5;
      else_7_else_1_equal_svs_st_6 <= else_7_else_1_equal_svs_st_5;
      else_7_equal_svs_st_6 <= else_7_equal_svs_st_5;
      max_sg1_lpi_dfm_3_st_6 <= max_sg1_lpi_dfm_3_st_5;
      if_7_equal_svs_st_6 <= if_7_equal_svs_st_5;
      max_conc_4_tmp_mut_21_sg1 <= max_conc_4_tmp_mut_20_sg1;
      else_7_if_conc_tmp_mut_21_sg1 <= else_7_if_conc_tmp_mut_20_sg1;
      max_conc_4_tmp_mut_29_sg1 <= max_conc_4_tmp_mut_28_sg1;
      else_7_if_conc_tmp_mut_29_sg1 <= else_7_if_conc_tmp_mut_28_sg1;
      max_conc_4_tmp_mut_37_sg1 <= max_conc_4_tmp_mut_36_sg1;
      else_7_if_conc_tmp_mut_37_sg1 <= else_7_if_conc_tmp_mut_36_sg1;
      max_conc_4_tmp_mut_45_sg1 <= max_conc_4_tmp_mut_44_sg1;
      else_7_if_conc_tmp_mut_45_sg1 <= else_7_if_conc_tmp_mut_44_sg1;
      max_conc_4_tmp_mut_53_sg1 <= max_conc_4_tmp_mut_52_sg1;
      else_7_if_conc_tmp_mut_53_sg1 <= else_7_if_conc_tmp_mut_52_sg1;
      max_conc_4_tmp_mut_61_sg1 <= max_conc_4_tmp_mut_60_sg1;
      else_7_if_conc_tmp_mut_61_sg1 <= else_7_if_conc_tmp_mut_60_sg1;
      max_conc_4_tmp_mut_69_sg1 <= max_conc_4_tmp_mut_68_sg1;
      else_7_if_conc_tmp_mut_69_sg1 <= else_7_if_conc_tmp_mut_68_sg1;
      max_conc_4_tmp_mut_77_sg1 <= max_conc_4_tmp_mut_76_sg1;
      else_7_if_conc_tmp_mut_77_sg1 <= else_7_if_conc_tmp_mut_76_sg1;
      max_conc_4_tmp_mut_13_sg1 <= max_conc_4_tmp_mut_12_sg1;
      else_7_if_conc_tmp_mut_13_sg1 <= else_7_if_conc_tmp_mut_12_sg1;
      else_7_if_div_9cyc_st_5 <= else_7_if_div_9cyc_st_4;
      delta_conc_1_tmp_mut_21_sg1 <= delta_conc_1_tmp_mut_20_sg1;
      else_7_if_1_conc_tmp_mut_21_sg1 <= else_7_if_1_conc_tmp_mut_20_sg1;
      delta_conc_1_tmp_mut_29_sg1 <= delta_conc_1_tmp_mut_28_sg1;
      else_7_if_1_conc_tmp_mut_29_sg1 <= else_7_if_1_conc_tmp_mut_28_sg1;
      delta_conc_1_tmp_mut_37_sg1 <= delta_conc_1_tmp_mut_36_sg1;
      else_7_if_1_conc_tmp_mut_37_sg1 <= else_7_if_1_conc_tmp_mut_36_sg1;
      delta_conc_1_tmp_mut_45_sg1 <= delta_conc_1_tmp_mut_44_sg1;
      else_7_if_1_conc_tmp_mut_45_sg1 <= else_7_if_1_conc_tmp_mut_44_sg1;
      delta_conc_1_tmp_mut_53_sg1 <= delta_conc_1_tmp_mut_52_sg1;
      else_7_if_1_conc_tmp_mut_53_sg1 <= else_7_if_1_conc_tmp_mut_52_sg1;
      delta_conc_1_tmp_mut_61_sg1 <= delta_conc_1_tmp_mut_60_sg1;
      else_7_if_1_conc_tmp_mut_61_sg1 <= else_7_if_1_conc_tmp_mut_60_sg1;
      delta_conc_1_tmp_mut_69_sg1 <= delta_conc_1_tmp_mut_68_sg1;
      else_7_if_1_conc_tmp_mut_69_sg1 <= else_7_if_1_conc_tmp_mut_68_sg1;
      delta_conc_1_tmp_mut_77_sg1 <= delta_conc_1_tmp_mut_76_sg1;
      else_7_if_1_conc_tmp_mut_77_sg1 <= else_7_if_1_conc_tmp_mut_76_sg1;
      delta_conc_1_tmp_mut_13_sg1 <= delta_conc_1_tmp_mut_12_sg1;
      else_7_if_1_conc_tmp_mut_13_sg1 <= else_7_if_1_conc_tmp_mut_12_sg1;
      else_7_if_1_div_9cyc_st_5 <= else_7_if_1_div_9cyc_st_4;
      delta_conc_2_tmp_mut_13_sg1 <= delta_conc_2_tmp_mut_12_sg1;
      else_7_else_1_if_conc_tmp_mut_13_sg1 <= else_7_else_1_if_conc_tmp_mut_12_sg1;
      delta_conc_2_tmp_mut_21_sg1 <= delta_conc_2_tmp_mut_20_sg1;
      else_7_else_1_if_conc_tmp_mut_21_sg1 <= else_7_else_1_if_conc_tmp_mut_20_sg1;
      delta_conc_2_tmp_mut_29_sg1 <= delta_conc_2_tmp_mut_28_sg1;
      else_7_else_1_if_conc_tmp_mut_29_sg1 <= else_7_else_1_if_conc_tmp_mut_28_sg1;
      delta_conc_2_tmp_mut_37_sg1 <= delta_conc_2_tmp_mut_36_sg1;
      else_7_else_1_if_conc_tmp_mut_37_sg1 <= else_7_else_1_if_conc_tmp_mut_36_sg1;
      delta_conc_2_tmp_mut_45_sg1 <= delta_conc_2_tmp_mut_44_sg1;
      else_7_else_1_if_conc_tmp_mut_45_sg1 <= else_7_else_1_if_conc_tmp_mut_44_sg1;
      delta_conc_2_tmp_mut_53_sg1 <= delta_conc_2_tmp_mut_52_sg1;
      else_7_else_1_if_conc_tmp_mut_53_sg1 <= else_7_else_1_if_conc_tmp_mut_52_sg1;
      delta_conc_2_tmp_mut_61_sg1 <= delta_conc_2_tmp_mut_60_sg1;
      else_7_else_1_if_conc_tmp_mut_61_sg1 <= else_7_else_1_if_conc_tmp_mut_60_sg1;
      delta_conc_2_tmp_mut_69_sg1 <= delta_conc_2_tmp_mut_68_sg1;
      else_7_else_1_if_conc_tmp_mut_69_sg1 <= else_7_else_1_if_conc_tmp_mut_68_sg1;
      delta_conc_2_tmp_mut_77_sg1 <= delta_conc_2_tmp_mut_76_sg1;
      else_7_else_1_if_conc_tmp_mut_77_sg1 <= else_7_else_1_if_conc_tmp_mut_76_sg1;
      else_7_else_1_if_div_9cyc_st_5 <= else_7_else_1_if_div_9cyc_st_4;
      delta_conc_3_tmp_mut_13_sg1 <= delta_conc_3_tmp_mut_12_sg1;
      else_7_else_1_else_conc_tmp_mut_13_sg1 <= else_7_else_1_else_conc_tmp_mut_12_sg1;
      delta_conc_3_tmp_mut_21_sg1 <= delta_conc_3_tmp_mut_20_sg1;
      else_7_else_1_else_conc_tmp_mut_21_sg1 <= else_7_else_1_else_conc_tmp_mut_20_sg1;
      delta_conc_3_tmp_mut_29_sg1 <= delta_conc_3_tmp_mut_28_sg1;
      else_7_else_1_else_conc_tmp_mut_29_sg1 <= else_7_else_1_else_conc_tmp_mut_28_sg1;
      delta_conc_3_tmp_mut_37_sg1 <= delta_conc_3_tmp_mut_36_sg1;
      else_7_else_1_else_conc_tmp_mut_37_sg1 <= else_7_else_1_else_conc_tmp_mut_36_sg1;
      delta_conc_3_tmp_mut_45_sg1 <= delta_conc_3_tmp_mut_44_sg1;
      else_7_else_1_else_conc_tmp_mut_45_sg1 <= else_7_else_1_else_conc_tmp_mut_44_sg1;
      delta_conc_3_tmp_mut_53_sg1 <= delta_conc_3_tmp_mut_52_sg1;
      else_7_else_1_else_conc_tmp_mut_53_sg1 <= else_7_else_1_else_conc_tmp_mut_52_sg1;
      delta_conc_3_tmp_mut_61_sg1 <= delta_conc_3_tmp_mut_60_sg1;
      else_7_else_1_else_conc_tmp_mut_61_sg1 <= else_7_else_1_else_conc_tmp_mut_60_sg1;
      delta_conc_3_tmp_mut_69_sg1 <= delta_conc_3_tmp_mut_68_sg1;
      else_7_else_1_else_conc_tmp_mut_69_sg1 <= else_7_else_1_else_conc_tmp_mut_68_sg1;
      delta_conc_3_tmp_mut_77_sg1 <= delta_conc_3_tmp_mut_76_sg1;
      else_7_else_1_else_conc_tmp_mut_77_sg1 <= else_7_else_1_else_conc_tmp_mut_76_sg1;
      else_7_else_1_else_div_9cyc_st_5 <= else_7_else_1_else_div_9cyc_st_4;
      else_7_else_1_equal_svs_st_5 <= else_7_else_1_equal_svs_st_4;
      else_7_equal_svs_st_5 <= else_7_equal_svs_st_4;
      max_sg1_lpi_dfm_3_st_5 <= max_sg1_lpi_dfm_3_st_4;
      if_7_equal_svs_st_5 <= if_7_equal_svs_st_4;
      max_conc_4_tmp_mut_20_sg1 <= max_conc_4_tmp_mut_19_sg1;
      else_7_if_conc_tmp_mut_20_sg1 <= else_7_if_conc_tmp_mut_19_sg1;
      max_conc_4_tmp_mut_28_sg1 <= max_conc_4_tmp_mut_27_sg1;
      else_7_if_conc_tmp_mut_28_sg1 <= else_7_if_conc_tmp_mut_27_sg1;
      max_conc_4_tmp_mut_36_sg1 <= max_conc_4_tmp_mut_35_sg1;
      else_7_if_conc_tmp_mut_36_sg1 <= else_7_if_conc_tmp_mut_35_sg1;
      max_conc_4_tmp_mut_44_sg1 <= max_conc_4_tmp_mut_43_sg1;
      else_7_if_conc_tmp_mut_44_sg1 <= else_7_if_conc_tmp_mut_43_sg1;
      max_conc_4_tmp_mut_52_sg1 <= max_conc_4_tmp_mut_51_sg1;
      else_7_if_conc_tmp_mut_52_sg1 <= else_7_if_conc_tmp_mut_51_sg1;
      max_conc_4_tmp_mut_60_sg1 <= max_conc_4_tmp_mut_59_sg1;
      else_7_if_conc_tmp_mut_60_sg1 <= else_7_if_conc_tmp_mut_59_sg1;
      max_conc_4_tmp_mut_68_sg1 <= max_conc_4_tmp_mut_67_sg1;
      else_7_if_conc_tmp_mut_68_sg1 <= else_7_if_conc_tmp_mut_67_sg1;
      max_conc_4_tmp_mut_76_sg1 <= max_conc_4_tmp_mut_75_sg1;
      else_7_if_conc_tmp_mut_76_sg1 <= else_7_if_conc_tmp_mut_75_sg1;
      max_conc_4_tmp_mut_12_sg1 <= max_conc_4_tmp_mut_11_sg1;
      else_7_if_conc_tmp_mut_12_sg1 <= else_7_if_conc_tmp_mut_11_sg1;
      else_7_if_div_9cyc_st_4 <= else_7_if_div_9cyc_st_3;
      delta_conc_1_tmp_mut_20_sg1 <= delta_conc_1_tmp_mut_19_sg1;
      else_7_if_1_conc_tmp_mut_20_sg1 <= else_7_if_1_conc_tmp_mut_19_sg1;
      delta_conc_1_tmp_mut_28_sg1 <= delta_conc_1_tmp_mut_27_sg1;
      else_7_if_1_conc_tmp_mut_28_sg1 <= else_7_if_1_conc_tmp_mut_27_sg1;
      delta_conc_1_tmp_mut_36_sg1 <= delta_conc_1_tmp_mut_35_sg1;
      else_7_if_1_conc_tmp_mut_36_sg1 <= else_7_if_1_conc_tmp_mut_35_sg1;
      delta_conc_1_tmp_mut_44_sg1 <= delta_conc_1_tmp_mut_43_sg1;
      else_7_if_1_conc_tmp_mut_44_sg1 <= else_7_if_1_conc_tmp_mut_43_sg1;
      delta_conc_1_tmp_mut_52_sg1 <= delta_conc_1_tmp_mut_51_sg1;
      else_7_if_1_conc_tmp_mut_52_sg1 <= else_7_if_1_conc_tmp_mut_51_sg1;
      delta_conc_1_tmp_mut_60_sg1 <= delta_conc_1_tmp_mut_59_sg1;
      else_7_if_1_conc_tmp_mut_60_sg1 <= else_7_if_1_conc_tmp_mut_59_sg1;
      delta_conc_1_tmp_mut_68_sg1 <= delta_conc_1_tmp_mut_67_sg1;
      else_7_if_1_conc_tmp_mut_68_sg1 <= else_7_if_1_conc_tmp_mut_67_sg1;
      delta_conc_1_tmp_mut_76_sg1 <= delta_conc_1_tmp_mut_75_sg1;
      else_7_if_1_conc_tmp_mut_76_sg1 <= else_7_if_1_conc_tmp_mut_75_sg1;
      delta_conc_1_tmp_mut_12_sg1 <= delta_conc_1_tmp_mut_11_sg1;
      else_7_if_1_conc_tmp_mut_12_sg1 <= else_7_if_1_conc_tmp_mut_11_sg1;
      else_7_if_1_div_9cyc_st_4 <= else_7_if_1_div_9cyc_st_3;
      delta_conc_2_tmp_mut_12_sg1 <= delta_conc_2_tmp_mut_11_sg1;
      else_7_else_1_if_conc_tmp_mut_12_sg1 <= else_7_else_1_if_conc_tmp_mut_11_sg1;
      delta_conc_2_tmp_mut_20_sg1 <= delta_conc_2_tmp_mut_19_sg1;
      else_7_else_1_if_conc_tmp_mut_20_sg1 <= else_7_else_1_if_conc_tmp_mut_19_sg1;
      delta_conc_2_tmp_mut_28_sg1 <= delta_conc_2_tmp_mut_27_sg1;
      else_7_else_1_if_conc_tmp_mut_28_sg1 <= else_7_else_1_if_conc_tmp_mut_27_sg1;
      delta_conc_2_tmp_mut_36_sg1 <= delta_conc_2_tmp_mut_35_sg1;
      else_7_else_1_if_conc_tmp_mut_36_sg1 <= else_7_else_1_if_conc_tmp_mut_35_sg1;
      delta_conc_2_tmp_mut_44_sg1 <= delta_conc_2_tmp_mut_43_sg1;
      else_7_else_1_if_conc_tmp_mut_44_sg1 <= else_7_else_1_if_conc_tmp_mut_43_sg1;
      delta_conc_2_tmp_mut_52_sg1 <= delta_conc_2_tmp_mut_51_sg1;
      else_7_else_1_if_conc_tmp_mut_52_sg1 <= else_7_else_1_if_conc_tmp_mut_51_sg1;
      delta_conc_2_tmp_mut_60_sg1 <= delta_conc_2_tmp_mut_59_sg1;
      else_7_else_1_if_conc_tmp_mut_60_sg1 <= else_7_else_1_if_conc_tmp_mut_59_sg1;
      delta_conc_2_tmp_mut_68_sg1 <= delta_conc_2_tmp_mut_67_sg1;
      else_7_else_1_if_conc_tmp_mut_68_sg1 <= else_7_else_1_if_conc_tmp_mut_67_sg1;
      delta_conc_2_tmp_mut_76_sg1 <= delta_conc_2_tmp_mut_75_sg1;
      else_7_else_1_if_conc_tmp_mut_76_sg1 <= else_7_else_1_if_conc_tmp_mut_75_sg1;
      else_7_else_1_if_div_9cyc_st_4 <= else_7_else_1_if_div_9cyc_st_3;
      delta_conc_3_tmp_mut_12_sg1 <= delta_conc_3_tmp_mut_11_sg1;
      else_7_else_1_else_conc_tmp_mut_12_sg1 <= else_7_else_1_else_conc_tmp_mut_11_sg1;
      delta_conc_3_tmp_mut_20_sg1 <= delta_conc_3_tmp_mut_19_sg1;
      else_7_else_1_else_conc_tmp_mut_20_sg1 <= else_7_else_1_else_conc_tmp_mut_19_sg1;
      delta_conc_3_tmp_mut_28_sg1 <= delta_conc_3_tmp_mut_27_sg1;
      else_7_else_1_else_conc_tmp_mut_28_sg1 <= else_7_else_1_else_conc_tmp_mut_27_sg1;
      delta_conc_3_tmp_mut_36_sg1 <= delta_conc_3_tmp_mut_35_sg1;
      else_7_else_1_else_conc_tmp_mut_36_sg1 <= else_7_else_1_else_conc_tmp_mut_35_sg1;
      delta_conc_3_tmp_mut_44_sg1 <= delta_conc_3_tmp_mut_43_sg1;
      else_7_else_1_else_conc_tmp_mut_44_sg1 <= else_7_else_1_else_conc_tmp_mut_43_sg1;
      delta_conc_3_tmp_mut_52_sg1 <= delta_conc_3_tmp_mut_51_sg1;
      else_7_else_1_else_conc_tmp_mut_52_sg1 <= else_7_else_1_else_conc_tmp_mut_51_sg1;
      delta_conc_3_tmp_mut_60_sg1 <= delta_conc_3_tmp_mut_59_sg1;
      else_7_else_1_else_conc_tmp_mut_60_sg1 <= else_7_else_1_else_conc_tmp_mut_59_sg1;
      delta_conc_3_tmp_mut_68_sg1 <= delta_conc_3_tmp_mut_67_sg1;
      else_7_else_1_else_conc_tmp_mut_68_sg1 <= else_7_else_1_else_conc_tmp_mut_67_sg1;
      delta_conc_3_tmp_mut_76_sg1 <= delta_conc_3_tmp_mut_75_sg1;
      else_7_else_1_else_conc_tmp_mut_76_sg1 <= else_7_else_1_else_conc_tmp_mut_75_sg1;
      else_7_else_1_else_div_9cyc_st_4 <= else_7_else_1_else_div_9cyc_st_3;
      else_7_else_1_equal_svs_st_4 <= else_7_else_1_equal_svs_st_3;
      else_7_equal_svs_st_4 <= else_7_equal_svs_st_3;
      max_sg1_lpi_dfm_3_st_4 <= max_sg1_lpi_dfm_3_st_3;
      if_7_equal_svs_st_4 <= if_7_equal_svs_st_3;
      max_conc_4_tmp_mut_19_sg1 <= max_conc_4_tmp_mut_18_sg1;
      else_7_if_conc_tmp_mut_19_sg1 <= else_7_if_conc_tmp_mut_18_sg1;
      max_conc_4_tmp_mut_27_sg1 <= max_conc_4_tmp_mut_26_sg1;
      else_7_if_conc_tmp_mut_27_sg1 <= else_7_if_conc_tmp_mut_26_sg1;
      max_conc_4_tmp_mut_35_sg1 <= max_conc_4_tmp_mut_34_sg1;
      else_7_if_conc_tmp_mut_35_sg1 <= else_7_if_conc_tmp_mut_34_sg1;
      max_conc_4_tmp_mut_43_sg1 <= max_conc_4_tmp_mut_42_sg1;
      else_7_if_conc_tmp_mut_43_sg1 <= else_7_if_conc_tmp_mut_42_sg1;
      max_conc_4_tmp_mut_51_sg1 <= max_conc_4_tmp_mut_50_sg1;
      else_7_if_conc_tmp_mut_51_sg1 <= else_7_if_conc_tmp_mut_50_sg1;
      max_conc_4_tmp_mut_59_sg1 <= max_conc_4_tmp_mut_58_sg1;
      else_7_if_conc_tmp_mut_59_sg1 <= else_7_if_conc_tmp_mut_58_sg1;
      max_conc_4_tmp_mut_67_sg1 <= max_conc_4_tmp_mut_66_sg1;
      else_7_if_conc_tmp_mut_67_sg1 <= else_7_if_conc_tmp_mut_66_sg1;
      max_conc_4_tmp_mut_75_sg1 <= max_conc_4_tmp_mut_74_sg1;
      else_7_if_conc_tmp_mut_75_sg1 <= else_7_if_conc_tmp_mut_74_sg1;
      max_conc_4_tmp_mut_11_sg1 <= max_conc_4_tmp_mut_10_sg1;
      else_7_if_conc_tmp_mut_11_sg1 <= else_7_if_conc_tmp_mut_10_sg1;
      else_7_if_div_9cyc_st_3 <= else_7_if_div_9cyc_st_2;
      delta_conc_1_tmp_mut_19_sg1 <= delta_conc_1_tmp_mut_18_sg1;
      else_7_if_1_conc_tmp_mut_19_sg1 <= else_7_if_1_conc_tmp_mut_18_sg1;
      delta_conc_1_tmp_mut_27_sg1 <= delta_conc_1_tmp_mut_26_sg1;
      else_7_if_1_conc_tmp_mut_27_sg1 <= else_7_if_1_conc_tmp_mut_26_sg1;
      delta_conc_1_tmp_mut_35_sg1 <= delta_conc_1_tmp_mut_34_sg1;
      else_7_if_1_conc_tmp_mut_35_sg1 <= else_7_if_1_conc_tmp_mut_34_sg1;
      delta_conc_1_tmp_mut_43_sg1 <= delta_conc_1_tmp_mut_42_sg1;
      else_7_if_1_conc_tmp_mut_43_sg1 <= else_7_if_1_conc_tmp_mut_42_sg1;
      delta_conc_1_tmp_mut_51_sg1 <= delta_conc_1_tmp_mut_50_sg1;
      else_7_if_1_conc_tmp_mut_51_sg1 <= else_7_if_1_conc_tmp_mut_50_sg1;
      delta_conc_1_tmp_mut_59_sg1 <= delta_conc_1_tmp_mut_58_sg1;
      else_7_if_1_conc_tmp_mut_59_sg1 <= else_7_if_1_conc_tmp_mut_58_sg1;
      delta_conc_1_tmp_mut_67_sg1 <= delta_conc_1_tmp_mut_66_sg1;
      else_7_if_1_conc_tmp_mut_67_sg1 <= else_7_if_1_conc_tmp_mut_66_sg1;
      delta_conc_1_tmp_mut_75_sg1 <= delta_conc_1_tmp_mut_74_sg1;
      else_7_if_1_conc_tmp_mut_75_sg1 <= else_7_if_1_conc_tmp_mut_74_sg1;
      delta_conc_1_tmp_mut_11_sg1 <= delta_conc_1_tmp_mut_10_sg1;
      else_7_if_1_conc_tmp_mut_11_sg1 <= else_7_if_1_conc_tmp_mut_10_sg1;
      else_7_if_1_div_9cyc_st_3 <= else_7_if_1_div_9cyc_st_2;
      delta_conc_2_tmp_mut_11_sg1 <= delta_conc_2_tmp_mut_10_sg1;
      else_7_else_1_if_conc_tmp_mut_11_sg1 <= else_7_else_1_if_conc_tmp_mut_10_sg1;
      delta_conc_2_tmp_mut_19_sg1 <= delta_conc_2_tmp_mut_18_sg1;
      else_7_else_1_if_conc_tmp_mut_19_sg1 <= else_7_else_1_if_conc_tmp_mut_18_sg1;
      delta_conc_2_tmp_mut_27_sg1 <= delta_conc_2_tmp_mut_26_sg1;
      else_7_else_1_if_conc_tmp_mut_27_sg1 <= else_7_else_1_if_conc_tmp_mut_26_sg1;
      delta_conc_2_tmp_mut_35_sg1 <= delta_conc_2_tmp_mut_34_sg1;
      else_7_else_1_if_conc_tmp_mut_35_sg1 <= else_7_else_1_if_conc_tmp_mut_34_sg1;
      delta_conc_2_tmp_mut_43_sg1 <= delta_conc_2_tmp_mut_42_sg1;
      else_7_else_1_if_conc_tmp_mut_43_sg1 <= else_7_else_1_if_conc_tmp_mut_42_sg1;
      delta_conc_2_tmp_mut_51_sg1 <= delta_conc_2_tmp_mut_50_sg1;
      else_7_else_1_if_conc_tmp_mut_51_sg1 <= else_7_else_1_if_conc_tmp_mut_50_sg1;
      delta_conc_2_tmp_mut_59_sg1 <= delta_conc_2_tmp_mut_58_sg1;
      else_7_else_1_if_conc_tmp_mut_59_sg1 <= else_7_else_1_if_conc_tmp_mut_58_sg1;
      delta_conc_2_tmp_mut_67_sg1 <= delta_conc_2_tmp_mut_66_sg1;
      else_7_else_1_if_conc_tmp_mut_67_sg1 <= else_7_else_1_if_conc_tmp_mut_66_sg1;
      delta_conc_2_tmp_mut_75_sg1 <= delta_conc_2_tmp_mut_74_sg1;
      else_7_else_1_if_conc_tmp_mut_75_sg1 <= else_7_else_1_if_conc_tmp_mut_74_sg1;
      else_7_else_1_if_div_9cyc_st_3 <= else_7_else_1_if_div_9cyc_st_2;
      delta_conc_3_tmp_mut_11_sg1 <= delta_conc_3_tmp_mut_10_sg1;
      else_7_else_1_else_conc_tmp_mut_11_sg1 <= else_7_else_1_else_conc_tmp_mut_10_sg1;
      delta_conc_3_tmp_mut_19_sg1 <= delta_conc_3_tmp_mut_18_sg1;
      else_7_else_1_else_conc_tmp_mut_19_sg1 <= else_7_else_1_else_conc_tmp_mut_18_sg1;
      delta_conc_3_tmp_mut_27_sg1 <= delta_conc_3_tmp_mut_26_sg1;
      else_7_else_1_else_conc_tmp_mut_27_sg1 <= else_7_else_1_else_conc_tmp_mut_26_sg1;
      delta_conc_3_tmp_mut_35_sg1 <= delta_conc_3_tmp_mut_34_sg1;
      else_7_else_1_else_conc_tmp_mut_35_sg1 <= else_7_else_1_else_conc_tmp_mut_34_sg1;
      delta_conc_3_tmp_mut_43_sg1 <= delta_conc_3_tmp_mut_42_sg1;
      else_7_else_1_else_conc_tmp_mut_43_sg1 <= else_7_else_1_else_conc_tmp_mut_42_sg1;
      delta_conc_3_tmp_mut_51_sg1 <= delta_conc_3_tmp_mut_50_sg1;
      else_7_else_1_else_conc_tmp_mut_51_sg1 <= else_7_else_1_else_conc_tmp_mut_50_sg1;
      delta_conc_3_tmp_mut_59_sg1 <= delta_conc_3_tmp_mut_58_sg1;
      else_7_else_1_else_conc_tmp_mut_59_sg1 <= else_7_else_1_else_conc_tmp_mut_58_sg1;
      delta_conc_3_tmp_mut_67_sg1 <= delta_conc_3_tmp_mut_66_sg1;
      else_7_else_1_else_conc_tmp_mut_67_sg1 <= else_7_else_1_else_conc_tmp_mut_66_sg1;
      delta_conc_3_tmp_mut_75_sg1 <= delta_conc_3_tmp_mut_74_sg1;
      else_7_else_1_else_conc_tmp_mut_75_sg1 <= else_7_else_1_else_conc_tmp_mut_74_sg1;
      else_7_else_1_else_div_9cyc_st_3 <= else_7_else_1_else_div_9cyc_st_2;
      else_7_else_1_equal_svs_st_3 <= else_7_else_1_equal_svs_st_2;
      else_7_equal_svs_st_3 <= else_7_equal_svs_st_2;
      max_sg1_lpi_dfm_3_st_3 <= max_sg1_lpi_dfm_3_st_2;
      if_7_equal_svs_st_3 <= if_7_equal_svs_st_2;
      max_conc_4_tmp_mut_18_sg1 <= max_conc_4_tmp_mut_17_sg1;
      else_7_if_conc_tmp_mut_18_sg1 <= else_7_if_conc_tmp_mut_17_sg1;
      max_conc_4_tmp_mut_26_sg1 <= max_conc_4_tmp_mut_25_sg1;
      else_7_if_conc_tmp_mut_26_sg1 <= else_7_if_conc_tmp_mut_25_sg1;
      max_conc_4_tmp_mut_34_sg1 <= max_conc_4_tmp_mut_33_sg1;
      else_7_if_conc_tmp_mut_34_sg1 <= else_7_if_conc_tmp_mut_33_sg1;
      max_conc_4_tmp_mut_42_sg1 <= max_conc_4_tmp_mut_41_sg1;
      else_7_if_conc_tmp_mut_42_sg1 <= else_7_if_conc_tmp_mut_41_sg1;
      max_conc_4_tmp_mut_50_sg1 <= max_conc_4_tmp_mut_49_sg1;
      else_7_if_conc_tmp_mut_50_sg1 <= else_7_if_conc_tmp_mut_49_sg1;
      max_conc_4_tmp_mut_58_sg1 <= max_conc_4_tmp_mut_57_sg1;
      else_7_if_conc_tmp_mut_58_sg1 <= else_7_if_conc_tmp_mut_57_sg1;
      max_conc_4_tmp_mut_66_sg1 <= max_conc_4_tmp_mut_65_sg1;
      else_7_if_conc_tmp_mut_66_sg1 <= else_7_if_conc_tmp_mut_65_sg1;
      max_conc_4_tmp_mut_74_sg1 <= max_conc_4_tmp_mut_73_sg1;
      else_7_if_conc_tmp_mut_74_sg1 <= else_7_if_conc_tmp_mut_73_sg1;
      max_conc_4_tmp_mut_10_sg1 <= max_conc_4_tmp_mut_9_sg1;
      else_7_if_conc_tmp_mut_10_sg1 <= else_7_if_conc_tmp_mut_9_sg1;
      else_7_if_div_9cyc_st_2 <= else_7_if_div_9cyc_st_1;
      delta_conc_1_tmp_mut_18_sg1 <= delta_conc_1_tmp_mut_17_sg1;
      else_7_if_1_conc_tmp_mut_18_sg1 <= else_7_if_1_conc_tmp_mut_17_sg1;
      delta_conc_1_tmp_mut_26_sg1 <= delta_conc_1_tmp_mut_25_sg1;
      else_7_if_1_conc_tmp_mut_26_sg1 <= else_7_if_1_conc_tmp_mut_25_sg1;
      delta_conc_1_tmp_mut_34_sg1 <= delta_conc_1_tmp_mut_33_sg1;
      else_7_if_1_conc_tmp_mut_34_sg1 <= else_7_if_1_conc_tmp_mut_33_sg1;
      delta_conc_1_tmp_mut_42_sg1 <= delta_conc_1_tmp_mut_41_sg1;
      else_7_if_1_conc_tmp_mut_42_sg1 <= else_7_if_1_conc_tmp_mut_41_sg1;
      delta_conc_1_tmp_mut_50_sg1 <= delta_conc_1_tmp_mut_49_sg1;
      else_7_if_1_conc_tmp_mut_50_sg1 <= else_7_if_1_conc_tmp_mut_49_sg1;
      delta_conc_1_tmp_mut_58_sg1 <= delta_conc_1_tmp_mut_57_sg1;
      else_7_if_1_conc_tmp_mut_58_sg1 <= else_7_if_1_conc_tmp_mut_57_sg1;
      delta_conc_1_tmp_mut_66_sg1 <= delta_conc_1_tmp_mut_65_sg1;
      else_7_if_1_conc_tmp_mut_66_sg1 <= else_7_if_1_conc_tmp_mut_65_sg1;
      delta_conc_1_tmp_mut_74_sg1 <= delta_conc_1_tmp_mut_73_sg1;
      else_7_if_1_conc_tmp_mut_74_sg1 <= else_7_if_1_conc_tmp_mut_73_sg1;
      delta_conc_1_tmp_mut_10_sg1 <= delta_conc_1_tmp_mut_9_sg1;
      else_7_if_1_conc_tmp_mut_10_sg1 <= else_7_if_1_conc_tmp_mut_9_sg1;
      else_7_if_1_div_9cyc_st_2 <= else_7_if_1_div_9cyc;
      delta_conc_2_tmp_mut_10_sg1 <= delta_conc_2_tmp_mut_9_sg1;
      else_7_else_1_if_conc_tmp_mut_10_sg1 <= else_7_else_1_if_conc_tmp_mut_9_sg1;
      delta_conc_2_tmp_mut_18_sg1 <= delta_conc_2_tmp_mut_17_sg1;
      else_7_else_1_if_conc_tmp_mut_18_sg1 <= else_7_else_1_if_conc_tmp_mut_17_sg1;
      delta_conc_2_tmp_mut_26_sg1 <= delta_conc_2_tmp_mut_25_sg1;
      else_7_else_1_if_conc_tmp_mut_26_sg1 <= else_7_else_1_if_conc_tmp_mut_25_sg1;
      delta_conc_2_tmp_mut_34_sg1 <= delta_conc_2_tmp_mut_33_sg1;
      else_7_else_1_if_conc_tmp_mut_34_sg1 <= else_7_else_1_if_conc_tmp_mut_33_sg1;
      delta_conc_2_tmp_mut_42_sg1 <= delta_conc_2_tmp_mut_41_sg1;
      else_7_else_1_if_conc_tmp_mut_42_sg1 <= else_7_else_1_if_conc_tmp_mut_41_sg1;
      delta_conc_2_tmp_mut_50_sg1 <= delta_conc_2_tmp_mut_49_sg1;
      else_7_else_1_if_conc_tmp_mut_50_sg1 <= else_7_else_1_if_conc_tmp_mut_49_sg1;
      delta_conc_2_tmp_mut_58_sg1 <= delta_conc_2_tmp_mut_57_sg1;
      else_7_else_1_if_conc_tmp_mut_58_sg1 <= else_7_else_1_if_conc_tmp_mut_57_sg1;
      delta_conc_2_tmp_mut_66_sg1 <= delta_conc_2_tmp_mut_65_sg1;
      else_7_else_1_if_conc_tmp_mut_66_sg1 <= else_7_else_1_if_conc_tmp_mut_65_sg1;
      delta_conc_2_tmp_mut_74_sg1 <= delta_conc_2_tmp_mut_73_sg1;
      else_7_else_1_if_conc_tmp_mut_74_sg1 <= else_7_else_1_if_conc_tmp_mut_73_sg1;
      else_7_else_1_if_div_9cyc_st_2 <= else_7_else_1_if_div_9cyc;
      delta_conc_3_tmp_mut_10_sg1 <= delta_conc_3_tmp_mut_9_sg1;
      else_7_else_1_else_conc_tmp_mut_10_sg1 <= else_7_else_1_else_conc_tmp_mut_9_sg1;
      delta_conc_3_tmp_mut_18_sg1 <= delta_conc_3_tmp_mut_17_sg1;
      else_7_else_1_else_conc_tmp_mut_18_sg1 <= else_7_else_1_else_conc_tmp_mut_17_sg1;
      delta_conc_3_tmp_mut_26_sg1 <= delta_conc_3_tmp_mut_25_sg1;
      else_7_else_1_else_conc_tmp_mut_26_sg1 <= else_7_else_1_else_conc_tmp_mut_25_sg1;
      delta_conc_3_tmp_mut_34_sg1 <= delta_conc_3_tmp_mut_33_sg1;
      else_7_else_1_else_conc_tmp_mut_34_sg1 <= else_7_else_1_else_conc_tmp_mut_33_sg1;
      delta_conc_3_tmp_mut_42_sg1 <= delta_conc_3_tmp_mut_41_sg1;
      else_7_else_1_else_conc_tmp_mut_42_sg1 <= else_7_else_1_else_conc_tmp_mut_41_sg1;
      delta_conc_3_tmp_mut_50_sg1 <= delta_conc_3_tmp_mut_49_sg1;
      else_7_else_1_else_conc_tmp_mut_50_sg1 <= else_7_else_1_else_conc_tmp_mut_49_sg1;
      delta_conc_3_tmp_mut_58_sg1 <= delta_conc_3_tmp_mut_57_sg1;
      else_7_else_1_else_conc_tmp_mut_58_sg1 <= else_7_else_1_else_conc_tmp_mut_57_sg1;
      delta_conc_3_tmp_mut_66_sg1 <= delta_conc_3_tmp_mut_65_sg1;
      else_7_else_1_else_conc_tmp_mut_66_sg1 <= else_7_else_1_else_conc_tmp_mut_65_sg1;
      delta_conc_3_tmp_mut_74_sg1 <= delta_conc_3_tmp_mut_73_sg1;
      else_7_else_1_else_conc_tmp_mut_74_sg1 <= else_7_else_1_else_conc_tmp_mut_73_sg1;
      else_7_else_1_else_div_9cyc_st_2 <= else_7_else_1_else_div_9cyc;
      else_7_else_1_equal_svs_st_2 <= else_7_else_1_equal_svs_1;
      else_7_equal_svs_st_2 <= else_7_equal_svs_st_1;
      max_sg1_lpi_dfm_3_st_2 <= max_sg1_lpi_dfm_3_st_1;
      if_7_equal_svs_st_2 <= if_7_equal_svs_st_1;
      max_conc_4_tmp_mut_17_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_17_sg1},
          or_4933_cse);
      else_7_if_conc_tmp_mut_17_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_17_sg1},
          or_4933_cse);
      max_conc_4_tmp_mut_25_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_25_sg1},
          or_4943_cse);
      else_7_if_conc_tmp_mut_25_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_25_sg1},
          or_4943_cse);
      max_conc_4_tmp_mut_33_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_33_sg1},
          or_4953_cse);
      else_7_if_conc_tmp_mut_33_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_33_sg1},
          or_4953_cse);
      max_conc_4_tmp_mut_41_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_41_sg1},
          or_4963_cse);
      else_7_if_conc_tmp_mut_41_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_41_sg1},
          or_4963_cse);
      max_conc_4_tmp_mut_49_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_49_sg1},
          or_4973_cse);
      else_7_if_conc_tmp_mut_49_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_49_sg1},
          or_4973_cse);
      max_conc_4_tmp_mut_57_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_57_sg1},
          or_4983_cse);
      else_7_if_conc_tmp_mut_57_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_57_sg1},
          or_4983_cse);
      max_conc_4_tmp_mut_65_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_65_sg1},
          or_4993_cse);
      else_7_if_conc_tmp_mut_65_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_65_sg1},
          or_4993_cse);
      max_conc_4_tmp_mut_73_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_73_sg1},
          or_5003_cse);
      else_7_if_conc_tmp_mut_73_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_73_sg1},
          or_5003_cse);
      max_conc_4_tmp_mut_9_sg1 <= MUX_v_16_2_2({mux1h_81_tmp , max_conc_4_tmp_mut_9_sg1},
          or_5013_cse);
      else_7_if_conc_tmp_mut_9_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_9_sg1},
          or_5013_cse);
      else_7_if_div_9cyc_st_1 <= MUX_v_4_2_2({else_7_if_acc_tmp , else_7_if_div_9cyc_st},
          and_9058_cse);
      delta_conc_1_tmp_mut_17_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_17_sg1},
          or_5023_cse);
      else_7_if_1_conc_tmp_mut_17_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_17_sg1}, or_5023_cse);
      delta_conc_1_tmp_mut_25_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_25_sg1},
          or_5033_cse);
      else_7_if_1_conc_tmp_mut_25_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_25_sg1}, or_5033_cse);
      delta_conc_1_tmp_mut_33_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_33_sg1},
          or_5043_cse);
      else_7_if_1_conc_tmp_mut_33_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_33_sg1}, or_5043_cse);
      delta_conc_1_tmp_mut_41_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_41_sg1},
          or_5053_cse);
      else_7_if_1_conc_tmp_mut_41_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_41_sg1}, or_5053_cse);
      delta_conc_1_tmp_mut_49_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_49_sg1},
          or_5063_cse);
      else_7_if_1_conc_tmp_mut_49_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_49_sg1}, or_5063_cse);
      delta_conc_1_tmp_mut_57_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_57_sg1},
          or_5073_cse);
      else_7_if_1_conc_tmp_mut_57_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_57_sg1}, or_5073_cse);
      delta_conc_1_tmp_mut_65_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_65_sg1},
          or_5083_cse);
      else_7_if_1_conc_tmp_mut_65_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_65_sg1}, or_5083_cse);
      delta_conc_1_tmp_mut_73_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_73_sg1},
          or_5093_cse);
      else_7_if_1_conc_tmp_mut_73_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_73_sg1}, or_5093_cse);
      delta_conc_1_tmp_mut_9_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_9_sg1},
          or_5103_cse);
      else_7_if_1_conc_tmp_mut_9_sg1 <= MUX_v_17_2_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_9_sg1}, or_5103_cse);
      delta_conc_2_tmp_mut_9_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_9_sg1},
          or_5114_cse);
      else_7_else_1_if_conc_tmp_mut_9_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_9_sg1}, or_5114_cse);
      delta_conc_2_tmp_mut_17_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_17_sg1},
          or_5126_cse);
      else_7_else_1_if_conc_tmp_mut_17_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_17_sg1}, or_5126_cse);
      delta_conc_2_tmp_mut_25_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_25_sg1},
          or_5138_cse);
      else_7_else_1_if_conc_tmp_mut_25_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_25_sg1}, or_5138_cse);
      delta_conc_2_tmp_mut_33_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_33_sg1},
          or_5150_cse);
      else_7_else_1_if_conc_tmp_mut_33_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_33_sg1}, or_5150_cse);
      delta_conc_2_tmp_mut_41_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_41_sg1},
          or_5162_cse);
      else_7_else_1_if_conc_tmp_mut_41_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_41_sg1}, or_5162_cse);
      delta_conc_2_tmp_mut_49_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_49_sg1},
          or_5174_cse);
      else_7_else_1_if_conc_tmp_mut_49_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_49_sg1}, or_5174_cse);
      delta_conc_2_tmp_mut_57_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_57_sg1},
          or_5186_cse);
      else_7_else_1_if_conc_tmp_mut_57_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_57_sg1}, or_5186_cse);
      delta_conc_2_tmp_mut_65_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_65_sg1},
          or_5198_cse);
      else_7_else_1_if_conc_tmp_mut_65_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_65_sg1}, or_5198_cse);
      delta_conc_2_tmp_mut_73_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_73_sg1},
          or_5210_cse);
      else_7_else_1_if_conc_tmp_mut_73_sg1 <= MUX_v_17_2_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_73_sg1}, or_5210_cse);
      delta_conc_3_tmp_mut_9_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_9_sg1},
          or_5222_cse);
      else_7_else_1_else_conc_tmp_mut_9_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_9_sg1}, or_5222_cse);
      delta_conc_3_tmp_mut_17_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_17_sg1},
          or_5234_cse);
      else_7_else_1_else_conc_tmp_mut_17_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_17_sg1}, or_5234_cse);
      delta_conc_3_tmp_mut_25_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_25_sg1},
          or_5246_cse);
      else_7_else_1_else_conc_tmp_mut_25_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_25_sg1}, or_5246_cse);
      delta_conc_3_tmp_mut_33_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_33_sg1},
          or_5258_cse);
      else_7_else_1_else_conc_tmp_mut_33_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_33_sg1}, or_5258_cse);
      delta_conc_3_tmp_mut_41_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_41_sg1},
          or_5270_cse);
      else_7_else_1_else_conc_tmp_mut_41_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_41_sg1}, or_5270_cse);
      delta_conc_3_tmp_mut_49_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_49_sg1},
          or_5282_cse);
      else_7_else_1_else_conc_tmp_mut_49_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_49_sg1}, or_5282_cse);
      delta_conc_3_tmp_mut_57_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_57_sg1},
          or_5294_cse);
      else_7_else_1_else_conc_tmp_mut_57_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_57_sg1}, or_5294_cse);
      delta_conc_3_tmp_mut_65_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_65_sg1},
          or_5306_cse);
      else_7_else_1_else_conc_tmp_mut_65_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_65_sg1}, or_5306_cse);
      delta_conc_3_tmp_mut_73_sg1 <= MUX_v_16_2_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_73_sg1},
          or_5318_cse);
      else_7_else_1_else_conc_tmp_mut_73_sg1 <= MUX_v_17_2_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_73_sg1}, or_5318_cse);
      else_7_equal_svs_st_1 <= else_7_equal_tmp;
      max_sg1_lpi_dfm_3_st_1 <= mux1h_81_tmp;
      if_7_equal_svs_st_1 <= if_7_equal_tmp;
      else_7_if_div_9cyc <= MUX_v_4_2_2({else_7_if_acc_tmp , else_7_if_div_9cyc},
          or_5325_cse);
      else_7_if_1_div_9cyc <= MUX_v_4_2_2({else_7_if_1_acc_tmp , else_7_if_1_div_9cyc},
          or_dcpl_856);
      else_7_else_1_if_div_9cyc <= MUX_v_4_2_2({else_7_else_1_if_acc_tmp , else_7_else_1_if_div_9cyc},
          or_dcpl_947 | (~ else_7_else_1_equal_tmp));
      else_7_else_1_else_div_9cyc <= MUX_v_4_2_2({else_7_else_1_else_acc_tmp , else_7_else_1_else_div_9cyc},
          or_dcpl_947 | else_7_else_1_equal_tmp);
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      main_stage_0_7 <= main_stage_0_6;
      main_stage_0_8 <= main_stage_0_7;
      main_stage_0_9 <= main_stage_0_8;
      main_stage_0_10 <= main_stage_0_9;
      else_7_if_div_9cyc_st <= MUX_v_4_2_2({else_7_if_acc_tmp , else_7_if_div_9cyc_st},
          or_5325_cse);
      slc_3_itm_8 <= slc_3_itm_7;
      else_7_and_5_itm_8 <= else_7_and_5_itm_7;
      unequal_tmp_8 <= unequal_tmp_7;
      slc_3_itm_7 <= slc_3_itm_6;
      else_7_and_5_itm_7 <= else_7_and_5_itm_6;
      unequal_tmp_7 <= unequal_tmp_6;
      slc_3_itm_6 <= slc_3_itm_5;
      else_7_and_5_itm_6 <= else_7_and_5_itm_5;
      unequal_tmp_6 <= unequal_tmp_5;
      slc_3_itm_5 <= slc_3_itm_4;
      else_7_and_5_itm_5 <= else_7_and_5_itm_4;
      unequal_tmp_5 <= unequal_tmp_4;
      slc_3_itm_4 <= slc_3_itm_3;
      else_7_and_5_itm_4 <= else_7_and_5_itm_3;
      unequal_tmp_4 <= unequal_tmp_3;
      slc_3_itm_3 <= slc_3_itm_2;
      else_7_and_5_itm_3 <= else_7_and_5_itm_2;
      unequal_tmp_3 <= unequal_tmp_2;
      slc_3_itm_2 <= slc_3_itm_1;
      else_7_and_5_itm_2 <= else_7_and_5_itm_1;
      unequal_tmp_2 <= unequal_tmp_1;
      slc_3_itm_1 <= readslicef_69_15_54(conv_s2u_138_69(69'b11001000110010010011001000001101100110010100010110111
          * conv_s2s_16_69(mux1h_81_tmp)));
      else_7_and_5_itm_1 <= else_7_else_1_equal_tmp & (~ else_7_equal_tmp);
      unequal_tmp_1 <= unequal_tmp;
      else_7_else_1_equal_svs_1 <= else_7_else_1_equal_tmp;
      reg_div_mgc_div_28_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_17_sg1
          , max_conc_4_tmp_mut_18_sg1 , max_conc_4_tmp_mut_19_sg1 , max_conc_4_tmp_mut_20_sg1
          , max_conc_4_tmp_mut_21_sg1 , max_conc_4_tmp_mut_22_sg1 , max_conc_4_tmp_mut_23_sg1
          , max_conc_4_tmp_mut_24_sg1}, {and_3159_cse , and_3165_cse , and_3172_cse
          , and_3180_cse , and_3189_cse , and_3199_cse , and_3209_cse , and_3221_cse
          , mux_106_cse});
      reg_div_mgc_div_28_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_17_sg1
          , else_7_if_conc_tmp_mut_18_sg1 , else_7_if_conc_tmp_mut_19_sg1 , else_7_if_conc_tmp_mut_20_sg1
          , else_7_if_conc_tmp_mut_21_sg1 , else_7_if_conc_tmp_mut_22_sg1 , else_7_if_conc_tmp_mut_23_sg1
          , else_7_if_conc_tmp_mut_24_sg1}, {and_3159_cse , and_3165_cse , and_3172_cse
          , and_3180_cse , and_3189_cse , and_3199_cse , and_3209_cse , and_3221_cse
          , mux_106_cse});
      reg_div_mgc_div_29_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_25_sg1
          , max_conc_4_tmp_mut_26_sg1 , max_conc_4_tmp_mut_27_sg1 , max_conc_4_tmp_mut_28_sg1
          , max_conc_4_tmp_mut_29_sg1 , max_conc_4_tmp_mut_30_sg1 , max_conc_4_tmp_mut_31_sg1
          , max_conc_4_tmp_mut_32_sg1}, {and_3299_cse , and_3305_cse , and_3312_cse
          , and_3320_cse , and_3329_cse , and_3339_cse , and_3349_cse , and_3361_cse
          , mux_135_cse});
      reg_div_mgc_div_29_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_25_sg1
          , else_7_if_conc_tmp_mut_26_sg1 , else_7_if_conc_tmp_mut_27_sg1 , else_7_if_conc_tmp_mut_28_sg1
          , else_7_if_conc_tmp_mut_29_sg1 , else_7_if_conc_tmp_mut_30_sg1 , else_7_if_conc_tmp_mut_31_sg1
          , else_7_if_conc_tmp_mut_32_sg1}, {and_3299_cse , and_3305_cse , and_3312_cse
          , and_3320_cse , and_3329_cse , and_3339_cse , and_3349_cse , and_3361_cse
          , mux_135_cse});
      reg_div_mgc_div_30_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_33_sg1
          , max_conc_4_tmp_mut_34_sg1 , max_conc_4_tmp_mut_35_sg1 , max_conc_4_tmp_mut_36_sg1
          , max_conc_4_tmp_mut_37_sg1 , max_conc_4_tmp_mut_38_sg1 , max_conc_4_tmp_mut_39_sg1
          , max_conc_4_tmp_mut_40_sg1}, {and_3439_cse , and_3445_cse , and_3452_cse
          , and_3460_cse , and_3469_cse , and_3479_cse , and_3489_cse , and_3501_cse
          , mux_164_cse});
      reg_div_mgc_div_30_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_33_sg1
          , else_7_if_conc_tmp_mut_34_sg1 , else_7_if_conc_tmp_mut_35_sg1 , else_7_if_conc_tmp_mut_36_sg1
          , else_7_if_conc_tmp_mut_37_sg1 , else_7_if_conc_tmp_mut_38_sg1 , else_7_if_conc_tmp_mut_39_sg1
          , else_7_if_conc_tmp_mut_40_sg1}, {and_3439_cse , and_3445_cse , and_3452_cse
          , and_3460_cse , and_3469_cse , and_3479_cse , and_3489_cse , and_3501_cse
          , mux_164_cse});
      reg_div_mgc_div_31_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_41_sg1
          , max_conc_4_tmp_mut_42_sg1 , max_conc_4_tmp_mut_43_sg1 , max_conc_4_tmp_mut_44_sg1
          , max_conc_4_tmp_mut_45_sg1 , max_conc_4_tmp_mut_46_sg1 , max_conc_4_tmp_mut_47_sg1
          , max_conc_4_tmp_mut_48_sg1}, {and_3579_cse , and_3585_cse , and_3592_cse
          , and_3600_cse , and_3609_cse , and_3619_cse , and_3629_cse , and_3641_cse
          , mux_194_cse});
      reg_div_mgc_div_31_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_41_sg1
          , else_7_if_conc_tmp_mut_42_sg1 , else_7_if_conc_tmp_mut_43_sg1 , else_7_if_conc_tmp_mut_44_sg1
          , else_7_if_conc_tmp_mut_45_sg1 , else_7_if_conc_tmp_mut_46_sg1 , else_7_if_conc_tmp_mut_47_sg1
          , else_7_if_conc_tmp_mut_48_sg1}, {and_3579_cse , and_3585_cse , and_3592_cse
          , and_3600_cse , and_3609_cse , and_3619_cse , and_3629_cse , and_3641_cse
          , mux_194_cse});
      reg_div_mgc_div_32_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_49_sg1
          , max_conc_4_tmp_mut_50_sg1 , max_conc_4_tmp_mut_51_sg1 , max_conc_4_tmp_mut_52_sg1
          , max_conc_4_tmp_mut_53_sg1 , max_conc_4_tmp_mut_54_sg1 , max_conc_4_tmp_mut_55_sg1
          , max_conc_4_tmp_mut_56_sg1}, {and_3719_cse , and_3725_cse , and_3732_cse
          , and_3740_cse , and_3749_cse , and_3759_cse , and_3769_cse , and_3781_cse
          , mux_224_cse});
      reg_div_mgc_div_32_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_49_sg1
          , else_7_if_conc_tmp_mut_50_sg1 , else_7_if_conc_tmp_mut_51_sg1 , else_7_if_conc_tmp_mut_52_sg1
          , else_7_if_conc_tmp_mut_53_sg1 , else_7_if_conc_tmp_mut_54_sg1 , else_7_if_conc_tmp_mut_55_sg1
          , else_7_if_conc_tmp_mut_56_sg1}, {and_3719_cse , and_3725_cse , and_3732_cse
          , and_3740_cse , and_3749_cse , and_3759_cse , and_3769_cse , and_3781_cse
          , mux_224_cse});
      reg_div_mgc_div_33_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_57_sg1
          , max_conc_4_tmp_mut_58_sg1 , max_conc_4_tmp_mut_59_sg1 , max_conc_4_tmp_mut_60_sg1
          , max_conc_4_tmp_mut_61_sg1 , max_conc_4_tmp_mut_62_sg1 , max_conc_4_tmp_mut_63_sg1
          , max_conc_4_tmp_mut_64_sg1}, {and_3859_cse , and_3865_cse , and_3872_cse
          , and_3880_cse , and_3889_cse , and_3899_cse , and_3909_cse , and_3921_cse
          , mux_253_cse});
      reg_div_mgc_div_33_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_57_sg1
          , else_7_if_conc_tmp_mut_58_sg1 , else_7_if_conc_tmp_mut_59_sg1 , else_7_if_conc_tmp_mut_60_sg1
          , else_7_if_conc_tmp_mut_61_sg1 , else_7_if_conc_tmp_mut_62_sg1 , else_7_if_conc_tmp_mut_63_sg1
          , else_7_if_conc_tmp_mut_64_sg1}, {and_3859_cse , and_3865_cse , and_3872_cse
          , and_3880_cse , and_3889_cse , and_3899_cse , and_3909_cse , and_3921_cse
          , mux_253_cse});
      reg_div_mgc_div_34_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_65_sg1
          , max_conc_4_tmp_mut_66_sg1 , max_conc_4_tmp_mut_67_sg1 , max_conc_4_tmp_mut_68_sg1
          , max_conc_4_tmp_mut_69_sg1 , max_conc_4_tmp_mut_70_sg1 , max_conc_4_tmp_mut_71_sg1
          , max_conc_4_tmp_mut_72_sg1}, {and_3999_cse , and_4005_cse , and_4012_cse
          , and_4020_cse , and_4029_cse , and_4039_cse , and_4049_cse , and_4061_cse
          , mux_282_cse});
      reg_div_mgc_div_34_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_65_sg1
          , else_7_if_conc_tmp_mut_66_sg1 , else_7_if_conc_tmp_mut_67_sg1 , else_7_if_conc_tmp_mut_68_sg1
          , else_7_if_conc_tmp_mut_69_sg1 , else_7_if_conc_tmp_mut_70_sg1 , else_7_if_conc_tmp_mut_71_sg1
          , else_7_if_conc_tmp_mut_72_sg1}, {and_3999_cse , and_4005_cse , and_4012_cse
          , and_4020_cse , and_4029_cse , and_4039_cse , and_4049_cse , and_4061_cse
          , mux_282_cse});
      reg_div_mgc_div_35_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_73_sg1
          , max_conc_4_tmp_mut_74_sg1 , max_conc_4_tmp_mut_75_sg1 , max_conc_4_tmp_mut_76_sg1
          , max_conc_4_tmp_mut_77_sg1 , max_conc_4_tmp_mut_78_sg1 , max_conc_4_tmp_mut_79_sg1
          , max_conc_4_tmp_mut_80_sg1}, {and_4139_cse , and_4145_cse , and_4152_cse
          , and_4160_cse , and_4169_cse , and_4179_cse , and_4189_cse , and_4201_cse
          , mux_312_cse});
      reg_div_mgc_div_35_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_73_sg1
          , else_7_if_conc_tmp_mut_74_sg1 , else_7_if_conc_tmp_mut_75_sg1 , else_7_if_conc_tmp_mut_76_sg1
          , else_7_if_conc_tmp_mut_77_sg1 , else_7_if_conc_tmp_mut_78_sg1 , else_7_if_conc_tmp_mut_79_sg1
          , else_7_if_conc_tmp_mut_80_sg1}, {and_4139_cse , and_4145_cse , and_4152_cse
          , and_4160_cse , and_4169_cse , and_4179_cse , and_4189_cse , and_4201_cse
          , mux_312_cse});
      reg_div_mgc_div_27_b_tmp <= MUX1HOT_v_16_9_2({mux1h_81_tmp , max_conc_4_tmp_mut_9_sg1
          , max_conc_4_tmp_mut_10_sg1 , max_conc_4_tmp_mut_11_sg1 , max_conc_4_tmp_mut_12_sg1
          , max_conc_4_tmp_mut_13_sg1 , max_conc_4_tmp_mut_14_sg1 , max_conc_4_tmp_mut_15_sg1
          , max_conc_4_tmp_mut_16_sg1}, {and_4279_cse , and_4285_cse , and_4291_cse
          , and_4298_cse , and_4307_cse , and_4317_cse , and_4327_cse , and_4339_cse
          , mux_345_cse});
      reg_div_mgc_div_27_a_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , else_7_if_conc_tmp_mut_9_sg1
          , else_7_if_conc_tmp_mut_10_sg1 , else_7_if_conc_tmp_mut_11_sg1 , else_7_if_conc_tmp_mut_12_sg1
          , else_7_if_conc_tmp_mut_13_sg1 , else_7_if_conc_tmp_mut_14_sg1 , else_7_if_conc_tmp_mut_15_sg1
          , else_7_if_conc_tmp_mut_16_sg1}, {and_4279_cse , and_4285_cse , and_4291_cse
          , and_4298_cse , and_4307_cse , and_4317_cse , and_4327_cse , and_4339_cse
          , mux_345_cse});
      reg_div_mgc_div_19_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_17_sg1
          , delta_conc_1_tmp_mut_18_sg1 , delta_conc_1_tmp_mut_19_sg1 , delta_conc_1_tmp_mut_20_sg1
          , delta_conc_1_tmp_mut_21_sg1 , delta_conc_1_tmp_mut_22_sg1 , delta_conc_1_tmp_mut_23_sg1
          , delta_conc_1_tmp_mut_24_sg1}, {and_4415_cse , and_4422_cse , and_4430_cse
          , and_4438_cse , and_4447_cse , and_4457_cse , and_4468_cse , and_4480_cse
          , and_4486_cse});
      reg_div_mgc_div_19_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_17_sg1 , else_7_if_1_conc_tmp_mut_18_sg1 , else_7_if_1_conc_tmp_mut_19_sg1
          , else_7_if_1_conc_tmp_mut_20_sg1 , else_7_if_1_conc_tmp_mut_21_sg1 , else_7_if_1_conc_tmp_mut_22_sg1
          , else_7_if_1_conc_tmp_mut_23_sg1 , else_7_if_1_conc_tmp_mut_24_sg1}, {and_4415_cse
          , and_4422_cse , and_4430_cse , and_4438_cse , and_4447_cse , and_4457_cse
          , and_4468_cse , and_4480_cse , and_4486_cse});
      reg_div_mgc_div_20_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_25_sg1
          , delta_conc_1_tmp_mut_26_sg1 , delta_conc_1_tmp_mut_27_sg1 , delta_conc_1_tmp_mut_28_sg1
          , delta_conc_1_tmp_mut_29_sg1 , delta_conc_1_tmp_mut_30_sg1 , delta_conc_1_tmp_mut_31_sg1
          , delta_conc_1_tmp_mut_32_sg1}, {and_4566_cse , and_4573_cse , and_4581_cse
          , and_4589_cse , and_4598_cse , and_4608_cse , and_4619_cse , and_4631_cse
          , and_4637_cse});
      reg_div_mgc_div_20_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_25_sg1 , else_7_if_1_conc_tmp_mut_26_sg1 , else_7_if_1_conc_tmp_mut_27_sg1
          , else_7_if_1_conc_tmp_mut_28_sg1 , else_7_if_1_conc_tmp_mut_29_sg1 , else_7_if_1_conc_tmp_mut_30_sg1
          , else_7_if_1_conc_tmp_mut_31_sg1 , else_7_if_1_conc_tmp_mut_32_sg1}, {and_4566_cse
          , and_4573_cse , and_4581_cse , and_4589_cse , and_4598_cse , and_4608_cse
          , and_4619_cse , and_4631_cse , and_4637_cse});
      reg_div_mgc_div_21_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_33_sg1
          , delta_conc_1_tmp_mut_34_sg1 , delta_conc_1_tmp_mut_35_sg1 , delta_conc_1_tmp_mut_36_sg1
          , delta_conc_1_tmp_mut_37_sg1 , delta_conc_1_tmp_mut_38_sg1 , delta_conc_1_tmp_mut_39_sg1
          , delta_conc_1_tmp_mut_40_sg1}, {and_4717_cse , and_4724_cse , and_4732_cse
          , and_4740_cse , and_4749_cse , and_4759_cse , and_4770_cse , and_4782_cse
          , and_4788_cse});
      reg_div_mgc_div_21_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_33_sg1 , else_7_if_1_conc_tmp_mut_34_sg1 , else_7_if_1_conc_tmp_mut_35_sg1
          , else_7_if_1_conc_tmp_mut_36_sg1 , else_7_if_1_conc_tmp_mut_37_sg1 , else_7_if_1_conc_tmp_mut_38_sg1
          , else_7_if_1_conc_tmp_mut_39_sg1 , else_7_if_1_conc_tmp_mut_40_sg1}, {and_4717_cse
          , and_4724_cse , and_4732_cse , and_4740_cse , and_4749_cse , and_4759_cse
          , and_4770_cse , and_4782_cse , and_4788_cse});
      reg_div_mgc_div_22_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_41_sg1
          , delta_conc_1_tmp_mut_42_sg1 , delta_conc_1_tmp_mut_43_sg1 , delta_conc_1_tmp_mut_44_sg1
          , delta_conc_1_tmp_mut_45_sg1 , delta_conc_1_tmp_mut_46_sg1 , delta_conc_1_tmp_mut_47_sg1
          , delta_conc_1_tmp_mut_48_sg1}, {and_4868_cse , and_4875_cse , and_4883_cse
          , and_4891_cse , and_4900_cse , and_4910_cse , and_4921_cse , and_4933_cse
          , and_4939_cse});
      reg_div_mgc_div_22_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_41_sg1 , else_7_if_1_conc_tmp_mut_42_sg1 , else_7_if_1_conc_tmp_mut_43_sg1
          , else_7_if_1_conc_tmp_mut_44_sg1 , else_7_if_1_conc_tmp_mut_45_sg1 , else_7_if_1_conc_tmp_mut_46_sg1
          , else_7_if_1_conc_tmp_mut_47_sg1 , else_7_if_1_conc_tmp_mut_48_sg1}, {and_4868_cse
          , and_4875_cse , and_4883_cse , and_4891_cse , and_4900_cse , and_4910_cse
          , and_4921_cse , and_4933_cse , and_4939_cse});
      reg_div_mgc_div_23_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_49_sg1
          , delta_conc_1_tmp_mut_50_sg1 , delta_conc_1_tmp_mut_51_sg1 , delta_conc_1_tmp_mut_52_sg1
          , delta_conc_1_tmp_mut_53_sg1 , delta_conc_1_tmp_mut_54_sg1 , delta_conc_1_tmp_mut_55_sg1
          , delta_conc_1_tmp_mut_56_sg1}, {and_5019_cse , and_5026_cse , and_5034_cse
          , and_5042_cse , and_5051_cse , and_5061_cse , and_5072_cse , and_5084_cse
          , and_5090_cse});
      reg_div_mgc_div_23_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_49_sg1 , else_7_if_1_conc_tmp_mut_50_sg1 , else_7_if_1_conc_tmp_mut_51_sg1
          , else_7_if_1_conc_tmp_mut_52_sg1 , else_7_if_1_conc_tmp_mut_53_sg1 , else_7_if_1_conc_tmp_mut_54_sg1
          , else_7_if_1_conc_tmp_mut_55_sg1 , else_7_if_1_conc_tmp_mut_56_sg1}, {and_5019_cse
          , and_5026_cse , and_5034_cse , and_5042_cse , and_5051_cse , and_5061_cse
          , and_5072_cse , and_5084_cse , and_5090_cse});
      reg_div_mgc_div_24_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_57_sg1
          , delta_conc_1_tmp_mut_58_sg1 , delta_conc_1_tmp_mut_59_sg1 , delta_conc_1_tmp_mut_60_sg1
          , delta_conc_1_tmp_mut_61_sg1 , delta_conc_1_tmp_mut_62_sg1 , delta_conc_1_tmp_mut_63_sg1
          , delta_conc_1_tmp_mut_64_sg1}, {and_5170_cse , and_5177_cse , and_5185_cse
          , and_5193_cse , and_5202_cse , and_5212_cse , and_5223_cse , and_5235_cse
          , and_5241_cse});
      reg_div_mgc_div_24_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_57_sg1 , else_7_if_1_conc_tmp_mut_58_sg1 , else_7_if_1_conc_tmp_mut_59_sg1
          , else_7_if_1_conc_tmp_mut_60_sg1 , else_7_if_1_conc_tmp_mut_61_sg1 , else_7_if_1_conc_tmp_mut_62_sg1
          , else_7_if_1_conc_tmp_mut_63_sg1 , else_7_if_1_conc_tmp_mut_64_sg1}, {and_5170_cse
          , and_5177_cse , and_5185_cse , and_5193_cse , and_5202_cse , and_5212_cse
          , and_5223_cse , and_5235_cse , and_5241_cse});
      reg_div_mgc_div_25_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_65_sg1
          , delta_conc_1_tmp_mut_66_sg1 , delta_conc_1_tmp_mut_67_sg1 , delta_conc_1_tmp_mut_68_sg1
          , delta_conc_1_tmp_mut_69_sg1 , delta_conc_1_tmp_mut_70_sg1 , delta_conc_1_tmp_mut_71_sg1
          , delta_conc_1_tmp_mut_72_sg1}, {and_5321_cse , and_5328_cse , and_5336_cse
          , and_5344_cse , and_5353_cse , and_5363_cse , and_5374_cse , and_5386_cse
          , and_5392_cse});
      reg_div_mgc_div_25_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_65_sg1 , else_7_if_1_conc_tmp_mut_66_sg1 , else_7_if_1_conc_tmp_mut_67_sg1
          , else_7_if_1_conc_tmp_mut_68_sg1 , else_7_if_1_conc_tmp_mut_69_sg1 , else_7_if_1_conc_tmp_mut_70_sg1
          , else_7_if_1_conc_tmp_mut_71_sg1 , else_7_if_1_conc_tmp_mut_72_sg1}, {and_5321_cse
          , and_5328_cse , and_5336_cse , and_5344_cse , and_5353_cse , and_5363_cse
          , and_5374_cse , and_5386_cse , and_5392_cse});
      reg_div_mgc_div_26_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_73_sg1
          , delta_conc_1_tmp_mut_74_sg1 , delta_conc_1_tmp_mut_75_sg1 , delta_conc_1_tmp_mut_76_sg1
          , delta_conc_1_tmp_mut_77_sg1 , delta_conc_1_tmp_mut_78_sg1 , delta_conc_1_tmp_mut_79_sg1
          , delta_conc_1_tmp_mut_80_sg1}, {and_5472_cse , and_5479_cse , and_5487_cse
          , and_5495_cse , and_5504_cse , and_5514_cse , and_5525_cse , and_5537_cse
          , and_5543_cse});
      reg_div_mgc_div_26_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1])
          , else_7_if_1_conc_tmp_mut_73_sg1 , else_7_if_1_conc_tmp_mut_74_sg1 , else_7_if_1_conc_tmp_mut_75_sg1
          , else_7_if_1_conc_tmp_mut_76_sg1 , else_7_if_1_conc_tmp_mut_77_sg1 , else_7_if_1_conc_tmp_mut_78_sg1
          , else_7_if_1_conc_tmp_mut_79_sg1 , else_7_if_1_conc_tmp_mut_80_sg1}, {and_5472_cse
          , and_5479_cse , and_5487_cse , and_5495_cse , and_5504_cse , and_5514_cse
          , and_5525_cse , and_5537_cse , and_5543_cse});
      reg_div_mgc_div_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_1_tmp_mut_9_sg1
          , delta_conc_1_tmp_mut_10_sg1 , delta_conc_1_tmp_mut_11_sg1 , delta_conc_1_tmp_mut_12_sg1
          , delta_conc_1_tmp_mut_13_sg1 , delta_conc_1_tmp_mut_14_sg1 , delta_conc_1_tmp_mut_15_sg1
          , delta_conc_1_tmp_mut_16_sg1}, {and_5623_cse , and_5630_cse , and_5638_cse
          , and_5645_cse , and_5652_cse , and_5659_cse , and_5666_cse , and_5674_cse
          , mux_483_cse});
      reg_div_mgc_div_a_tmp <= MUX1HOT_v_17_9_2({(else_7_if_1_acc_1_itm[17:1]) ,
          else_7_if_1_conc_tmp_mut_9_sg1 , else_7_if_1_conc_tmp_mut_10_sg1 , else_7_if_1_conc_tmp_mut_11_sg1
          , else_7_if_1_conc_tmp_mut_12_sg1 , else_7_if_1_conc_tmp_mut_13_sg1 , else_7_if_1_conc_tmp_mut_14_sg1
          , else_7_if_1_conc_tmp_mut_15_sg1 , else_7_if_1_conc_tmp_mut_16_sg1}, {and_5623_cse
          , and_5630_cse , and_5638_cse , and_5645_cse , and_5652_cse , and_5659_cse
          , and_5666_cse , and_5674_cse , mux_483_cse});
      reg_div_mgc_div_10_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_9_sg1
          , delta_conc_2_tmp_mut_10_sg1 , delta_conc_2_tmp_mut_11_sg1 , delta_conc_2_tmp_mut_12_sg1
          , delta_conc_2_tmp_mut_13_sg1 , delta_conc_2_tmp_mut_14_sg1 , delta_conc_2_tmp_mut_15_sg1
          , delta_conc_2_tmp_mut_16_sg1}, {and_5737_cse , and_5745_cse , and_5754_cse
          , and_5763_cse , and_5773_cse , and_5784_cse , and_5796_cse , and_5809_cse
          , mux_514_cse});
      reg_div_mgc_div_10_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_9_sg1 , else_7_else_1_if_conc_tmp_mut_10_sg1
          , else_7_else_1_if_conc_tmp_mut_11_sg1 , else_7_else_1_if_conc_tmp_mut_12_sg1
          , else_7_else_1_if_conc_tmp_mut_13_sg1 , else_7_else_1_if_conc_tmp_mut_14_sg1
          , else_7_else_1_if_conc_tmp_mut_15_sg1 , else_7_else_1_if_conc_tmp_mut_16_sg1},
          {and_5737_cse , and_5745_cse , and_5754_cse , and_5763_cse , and_5773_cse
          , and_5784_cse , and_5796_cse , and_5809_cse , mux_514_cse});
      reg_div_mgc_div_11_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_17_sg1
          , delta_conc_2_tmp_mut_18_sg1 , delta_conc_2_tmp_mut_19_sg1 , delta_conc_2_tmp_mut_20_sg1
          , delta_conc_2_tmp_mut_21_sg1 , delta_conc_2_tmp_mut_22_sg1 , delta_conc_2_tmp_mut_23_sg1
          , delta_conc_2_tmp_mut_24_sg1}, {and_5904_cse , and_5912_cse , and_5921_cse
          , and_5930_cse , and_5940_cse , and_5951_cse , and_5963_cse , and_5976_cse
          , mux_526_cse});
      reg_div_mgc_div_11_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_17_sg1 , else_7_else_1_if_conc_tmp_mut_18_sg1
          , else_7_else_1_if_conc_tmp_mut_19_sg1 , else_7_else_1_if_conc_tmp_mut_20_sg1
          , else_7_else_1_if_conc_tmp_mut_21_sg1 , else_7_else_1_if_conc_tmp_mut_22_sg1
          , else_7_else_1_if_conc_tmp_mut_23_sg1 , else_7_else_1_if_conc_tmp_mut_24_sg1},
          {and_5904_cse , and_5912_cse , and_5921_cse , and_5930_cse , and_5940_cse
          , and_5951_cse , and_5963_cse , and_5976_cse , mux_526_cse});
      reg_div_mgc_div_12_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_25_sg1
          , delta_conc_2_tmp_mut_26_sg1 , delta_conc_2_tmp_mut_27_sg1 , delta_conc_2_tmp_mut_28_sg1
          , delta_conc_2_tmp_mut_29_sg1 , delta_conc_2_tmp_mut_30_sg1 , delta_conc_2_tmp_mut_31_sg1
          , delta_conc_2_tmp_mut_32_sg1}, {and_6071_cse , and_6079_cse , and_6088_cse
          , and_6097_cse , and_6107_cse , and_6118_cse , and_6130_cse , and_6143_cse
          , mux_538_cse});
      reg_div_mgc_div_12_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_25_sg1 , else_7_else_1_if_conc_tmp_mut_26_sg1
          , else_7_else_1_if_conc_tmp_mut_27_sg1 , else_7_else_1_if_conc_tmp_mut_28_sg1
          , else_7_else_1_if_conc_tmp_mut_29_sg1 , else_7_else_1_if_conc_tmp_mut_30_sg1
          , else_7_else_1_if_conc_tmp_mut_31_sg1 , else_7_else_1_if_conc_tmp_mut_32_sg1},
          {and_6071_cse , and_6079_cse , and_6088_cse , and_6097_cse , and_6107_cse
          , and_6118_cse , and_6130_cse , and_6143_cse , mux_538_cse});
      reg_div_mgc_div_13_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_33_sg1
          , delta_conc_2_tmp_mut_34_sg1 , delta_conc_2_tmp_mut_35_sg1 , delta_conc_2_tmp_mut_36_sg1
          , delta_conc_2_tmp_mut_37_sg1 , delta_conc_2_tmp_mut_38_sg1 , delta_conc_2_tmp_mut_39_sg1
          , delta_conc_2_tmp_mut_40_sg1}, {and_6238_cse , and_6246_cse , and_6255_cse
          , and_6264_cse , and_6274_cse , and_6285_cse , and_6297_cse , and_6310_cse
          , mux_550_cse});
      reg_div_mgc_div_13_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_33_sg1 , else_7_else_1_if_conc_tmp_mut_34_sg1
          , else_7_else_1_if_conc_tmp_mut_35_sg1 , else_7_else_1_if_conc_tmp_mut_36_sg1
          , else_7_else_1_if_conc_tmp_mut_37_sg1 , else_7_else_1_if_conc_tmp_mut_38_sg1
          , else_7_else_1_if_conc_tmp_mut_39_sg1 , else_7_else_1_if_conc_tmp_mut_40_sg1},
          {and_6238_cse , and_6246_cse , and_6255_cse , and_6264_cse , and_6274_cse
          , and_6285_cse , and_6297_cse , and_6310_cse , mux_550_cse});
      reg_div_mgc_div_14_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_41_sg1
          , delta_conc_2_tmp_mut_42_sg1 , delta_conc_2_tmp_mut_43_sg1 , delta_conc_2_tmp_mut_44_sg1
          , delta_conc_2_tmp_mut_45_sg1 , delta_conc_2_tmp_mut_46_sg1 , delta_conc_2_tmp_mut_47_sg1
          , delta_conc_2_tmp_mut_48_sg1}, {and_6405_cse , and_6413_cse , and_6422_cse
          , and_6431_cse , and_6441_cse , and_6452_cse , and_6464_cse , and_6477_cse
          , mux_562_cse});
      reg_div_mgc_div_14_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_41_sg1 , else_7_else_1_if_conc_tmp_mut_42_sg1
          , else_7_else_1_if_conc_tmp_mut_43_sg1 , else_7_else_1_if_conc_tmp_mut_44_sg1
          , else_7_else_1_if_conc_tmp_mut_45_sg1 , else_7_else_1_if_conc_tmp_mut_46_sg1
          , else_7_else_1_if_conc_tmp_mut_47_sg1 , else_7_else_1_if_conc_tmp_mut_48_sg1},
          {and_6405_cse , and_6413_cse , and_6422_cse , and_6431_cse , and_6441_cse
          , and_6452_cse , and_6464_cse , and_6477_cse , mux_562_cse});
      reg_div_mgc_div_15_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_49_sg1
          , delta_conc_2_tmp_mut_50_sg1 , delta_conc_2_tmp_mut_51_sg1 , delta_conc_2_tmp_mut_52_sg1
          , delta_conc_2_tmp_mut_53_sg1 , delta_conc_2_tmp_mut_54_sg1 , delta_conc_2_tmp_mut_55_sg1
          , delta_conc_2_tmp_mut_56_sg1}, {and_6572_cse , and_6580_cse , and_6589_cse
          , and_6598_cse , and_6608_cse , and_6619_cse , and_6631_cse , and_6644_cse
          , mux_574_cse});
      reg_div_mgc_div_15_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_49_sg1 , else_7_else_1_if_conc_tmp_mut_50_sg1
          , else_7_else_1_if_conc_tmp_mut_51_sg1 , else_7_else_1_if_conc_tmp_mut_52_sg1
          , else_7_else_1_if_conc_tmp_mut_53_sg1 , else_7_else_1_if_conc_tmp_mut_54_sg1
          , else_7_else_1_if_conc_tmp_mut_55_sg1 , else_7_else_1_if_conc_tmp_mut_56_sg1},
          {and_6572_cse , and_6580_cse , and_6589_cse , and_6598_cse , and_6608_cse
          , and_6619_cse , and_6631_cse , and_6644_cse , mux_574_cse});
      reg_div_mgc_div_16_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_57_sg1
          , delta_conc_2_tmp_mut_58_sg1 , delta_conc_2_tmp_mut_59_sg1 , delta_conc_2_tmp_mut_60_sg1
          , delta_conc_2_tmp_mut_61_sg1 , delta_conc_2_tmp_mut_62_sg1 , delta_conc_2_tmp_mut_63_sg1
          , delta_conc_2_tmp_mut_64_sg1}, {and_6739_cse , and_6747_cse , and_6756_cse
          , and_6765_cse , and_6775_cse , and_6786_cse , and_6798_cse , and_6811_cse
          , mux_586_cse});
      reg_div_mgc_div_16_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_57_sg1 , else_7_else_1_if_conc_tmp_mut_58_sg1
          , else_7_else_1_if_conc_tmp_mut_59_sg1 , else_7_else_1_if_conc_tmp_mut_60_sg1
          , else_7_else_1_if_conc_tmp_mut_61_sg1 , else_7_else_1_if_conc_tmp_mut_62_sg1
          , else_7_else_1_if_conc_tmp_mut_63_sg1 , else_7_else_1_if_conc_tmp_mut_64_sg1},
          {and_6739_cse , and_6747_cse , and_6756_cse , and_6765_cse , and_6775_cse
          , and_6786_cse , and_6798_cse , and_6811_cse , mux_586_cse});
      reg_div_mgc_div_17_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_65_sg1
          , delta_conc_2_tmp_mut_66_sg1 , delta_conc_2_tmp_mut_67_sg1 , delta_conc_2_tmp_mut_68_sg1
          , delta_conc_2_tmp_mut_69_sg1 , delta_conc_2_tmp_mut_70_sg1 , delta_conc_2_tmp_mut_71_sg1
          , delta_conc_2_tmp_mut_72_sg1}, {and_6906_cse , and_6914_cse , and_6923_cse
          , and_6932_cse , and_6942_cse , and_6953_cse , and_6965_cse , and_6978_cse
          , mux_598_cse});
      reg_div_mgc_div_17_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_65_sg1 , else_7_else_1_if_conc_tmp_mut_66_sg1
          , else_7_else_1_if_conc_tmp_mut_67_sg1 , else_7_else_1_if_conc_tmp_mut_68_sg1
          , else_7_else_1_if_conc_tmp_mut_69_sg1 , else_7_else_1_if_conc_tmp_mut_70_sg1
          , else_7_else_1_if_conc_tmp_mut_71_sg1 , else_7_else_1_if_conc_tmp_mut_72_sg1},
          {and_6906_cse , and_6914_cse , and_6923_cse , and_6932_cse , and_6942_cse
          , and_6953_cse , and_6965_cse , and_6978_cse , mux_598_cse});
      reg_div_mgc_div_18_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_2_tmp_mut_73_sg1
          , delta_conc_2_tmp_mut_74_sg1 , delta_conc_2_tmp_mut_75_sg1 , delta_conc_2_tmp_mut_76_sg1
          , delta_conc_2_tmp_mut_77_sg1 , delta_conc_2_tmp_mut_78_sg1 , delta_conc_2_tmp_mut_79_sg1
          , delta_conc_2_tmp_mut_80_sg1}, {and_7073_cse , and_7081_cse , and_7090_cse
          , and_7099_cse , and_7108_cse , and_7116_cse , and_7124_cse , and_7132_cse
          , mux_628_cse});
      reg_div_mgc_div_18_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_if_acc_2_itm[17:1])
          , else_7_else_1_if_conc_tmp_mut_73_sg1 , else_7_else_1_if_conc_tmp_mut_74_sg1
          , else_7_else_1_if_conc_tmp_mut_75_sg1 , else_7_else_1_if_conc_tmp_mut_76_sg1
          , else_7_else_1_if_conc_tmp_mut_77_sg1 , else_7_else_1_if_conc_tmp_mut_78_sg1
          , else_7_else_1_if_conc_tmp_mut_79_sg1 , else_7_else_1_if_conc_tmp_mut_80_sg1},
          {and_7073_cse , and_7081_cse , and_7090_cse , and_7099_cse , and_7108_cse
          , and_7116_cse , and_7124_cse , and_7132_cse , mux_628_cse});
      reg_div_mgc_div_1_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_9_sg1
          , delta_conc_3_tmp_mut_10_sg1 , delta_conc_3_tmp_mut_11_sg1 , delta_conc_3_tmp_mut_12_sg1
          , delta_conc_3_tmp_mut_13_sg1 , delta_conc_3_tmp_mut_14_sg1 , delta_conc_3_tmp_mut_15_sg1
          , delta_conc_3_tmp_mut_16_sg1}, {and_7204_cse , and_7212_cse , and_7221_cse
          , and_7231_cse , and_7242_cse , and_7254_cse , and_7267_cse , and_7281_cse
          , and_7288_cse});
      reg_div_mgc_div_1_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_9_sg1 , else_7_else_1_else_conc_tmp_mut_10_sg1
          , else_7_else_1_else_conc_tmp_mut_11_sg1 , else_7_else_1_else_conc_tmp_mut_12_sg1
          , else_7_else_1_else_conc_tmp_mut_13_sg1 , else_7_else_1_else_conc_tmp_mut_14_sg1
          , else_7_else_1_else_conc_tmp_mut_15_sg1 , else_7_else_1_else_conc_tmp_mut_16_sg1},
          {and_7204_cse , and_7212_cse , and_7221_cse , and_7231_cse , and_7242_cse
          , and_7254_cse , and_7267_cse , and_7281_cse , and_7288_cse});
      reg_div_mgc_div_2_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_17_sg1
          , delta_conc_3_tmp_mut_18_sg1 , delta_conc_3_tmp_mut_19_sg1 , delta_conc_3_tmp_mut_20_sg1
          , delta_conc_3_tmp_mut_21_sg1 , delta_conc_3_tmp_mut_22_sg1 , delta_conc_3_tmp_mut_23_sg1
          , delta_conc_3_tmp_mut_24_sg1}, {and_7383_cse , and_7391_cse , and_7400_cse
          , and_7410_cse , and_7421_cse , and_7433_cse , and_7446_cse , and_7460_cse
          , and_7467_cse});
      reg_div_mgc_div_2_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_17_sg1 , else_7_else_1_else_conc_tmp_mut_18_sg1
          , else_7_else_1_else_conc_tmp_mut_19_sg1 , else_7_else_1_else_conc_tmp_mut_20_sg1
          , else_7_else_1_else_conc_tmp_mut_21_sg1 , else_7_else_1_else_conc_tmp_mut_22_sg1
          , else_7_else_1_else_conc_tmp_mut_23_sg1 , else_7_else_1_else_conc_tmp_mut_24_sg1},
          {and_7383_cse , and_7391_cse , and_7400_cse , and_7410_cse , and_7421_cse
          , and_7433_cse , and_7446_cse , and_7460_cse , and_7467_cse});
      reg_div_mgc_div_3_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_25_sg1
          , delta_conc_3_tmp_mut_26_sg1 , delta_conc_3_tmp_mut_27_sg1 , delta_conc_3_tmp_mut_28_sg1
          , delta_conc_3_tmp_mut_29_sg1 , delta_conc_3_tmp_mut_30_sg1 , delta_conc_3_tmp_mut_31_sg1
          , delta_conc_3_tmp_mut_32_sg1}, {and_7562_cse , and_7570_cse , and_7579_cse
          , and_7589_cse , and_7600_cse , and_7612_cse , and_7625_cse , and_7639_cse
          , and_7646_cse});
      reg_div_mgc_div_3_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_25_sg1 , else_7_else_1_else_conc_tmp_mut_26_sg1
          , else_7_else_1_else_conc_tmp_mut_27_sg1 , else_7_else_1_else_conc_tmp_mut_28_sg1
          , else_7_else_1_else_conc_tmp_mut_29_sg1 , else_7_else_1_else_conc_tmp_mut_30_sg1
          , else_7_else_1_else_conc_tmp_mut_31_sg1 , else_7_else_1_else_conc_tmp_mut_32_sg1},
          {and_7562_cse , and_7570_cse , and_7579_cse , and_7589_cse , and_7600_cse
          , and_7612_cse , and_7625_cse , and_7639_cse , and_7646_cse});
      reg_div_mgc_div_4_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_33_sg1
          , delta_conc_3_tmp_mut_34_sg1 , delta_conc_3_tmp_mut_35_sg1 , delta_conc_3_tmp_mut_36_sg1
          , delta_conc_3_tmp_mut_37_sg1 , delta_conc_3_tmp_mut_38_sg1 , delta_conc_3_tmp_mut_39_sg1
          , delta_conc_3_tmp_mut_40_sg1}, {and_7741_cse , and_7749_cse , and_7758_cse
          , and_7768_cse , and_7779_cse , and_7791_cse , and_7804_cse , and_7818_cse
          , and_7825_cse});
      reg_div_mgc_div_4_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_33_sg1 , else_7_else_1_else_conc_tmp_mut_34_sg1
          , else_7_else_1_else_conc_tmp_mut_35_sg1 , else_7_else_1_else_conc_tmp_mut_36_sg1
          , else_7_else_1_else_conc_tmp_mut_37_sg1 , else_7_else_1_else_conc_tmp_mut_38_sg1
          , else_7_else_1_else_conc_tmp_mut_39_sg1 , else_7_else_1_else_conc_tmp_mut_40_sg1},
          {and_7741_cse , and_7749_cse , and_7758_cse , and_7768_cse , and_7779_cse
          , and_7791_cse , and_7804_cse , and_7818_cse , and_7825_cse});
      reg_div_mgc_div_5_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_41_sg1
          , delta_conc_3_tmp_mut_42_sg1 , delta_conc_3_tmp_mut_43_sg1 , delta_conc_3_tmp_mut_44_sg1
          , delta_conc_3_tmp_mut_45_sg1 , delta_conc_3_tmp_mut_46_sg1 , delta_conc_3_tmp_mut_47_sg1
          , delta_conc_3_tmp_mut_48_sg1}, {and_7920_cse , and_7928_cse , and_7937_cse
          , and_7947_cse , and_7958_cse , and_7970_cse , and_7983_cse , and_7997_cse
          , and_8004_cse});
      reg_div_mgc_div_5_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_41_sg1 , else_7_else_1_else_conc_tmp_mut_42_sg1
          , else_7_else_1_else_conc_tmp_mut_43_sg1 , else_7_else_1_else_conc_tmp_mut_44_sg1
          , else_7_else_1_else_conc_tmp_mut_45_sg1 , else_7_else_1_else_conc_tmp_mut_46_sg1
          , else_7_else_1_else_conc_tmp_mut_47_sg1 , else_7_else_1_else_conc_tmp_mut_48_sg1},
          {and_7920_cse , and_7928_cse , and_7937_cse , and_7947_cse , and_7958_cse
          , and_7970_cse , and_7983_cse , and_7997_cse , and_8004_cse});
      reg_div_mgc_div_6_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_49_sg1
          , delta_conc_3_tmp_mut_50_sg1 , delta_conc_3_tmp_mut_51_sg1 , delta_conc_3_tmp_mut_52_sg1
          , delta_conc_3_tmp_mut_53_sg1 , delta_conc_3_tmp_mut_54_sg1 , delta_conc_3_tmp_mut_55_sg1
          , delta_conc_3_tmp_mut_56_sg1}, {and_8099_cse , and_8107_cse , and_8116_cse
          , and_8126_cse , and_8137_cse , and_8149_cse , and_8162_cse , and_8176_cse
          , and_8183_cse});
      reg_div_mgc_div_6_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_49_sg1 , else_7_else_1_else_conc_tmp_mut_50_sg1
          , else_7_else_1_else_conc_tmp_mut_51_sg1 , else_7_else_1_else_conc_tmp_mut_52_sg1
          , else_7_else_1_else_conc_tmp_mut_53_sg1 , else_7_else_1_else_conc_tmp_mut_54_sg1
          , else_7_else_1_else_conc_tmp_mut_55_sg1 , else_7_else_1_else_conc_tmp_mut_56_sg1},
          {and_8099_cse , and_8107_cse , and_8116_cse , and_8126_cse , and_8137_cse
          , and_8149_cse , and_8162_cse , and_8176_cse , and_8183_cse});
      reg_div_mgc_div_7_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_57_sg1
          , delta_conc_3_tmp_mut_58_sg1 , delta_conc_3_tmp_mut_59_sg1 , delta_conc_3_tmp_mut_60_sg1
          , delta_conc_3_tmp_mut_61_sg1 , delta_conc_3_tmp_mut_62_sg1 , delta_conc_3_tmp_mut_63_sg1
          , delta_conc_3_tmp_mut_64_sg1}, {and_8278_cse , and_8286_cse , and_8295_cse
          , and_8305_cse , and_8316_cse , and_8328_cse , and_8341_cse , and_8355_cse
          , and_8362_cse});
      reg_div_mgc_div_7_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_57_sg1 , else_7_else_1_else_conc_tmp_mut_58_sg1
          , else_7_else_1_else_conc_tmp_mut_59_sg1 , else_7_else_1_else_conc_tmp_mut_60_sg1
          , else_7_else_1_else_conc_tmp_mut_61_sg1 , else_7_else_1_else_conc_tmp_mut_62_sg1
          , else_7_else_1_else_conc_tmp_mut_63_sg1 , else_7_else_1_else_conc_tmp_mut_64_sg1},
          {and_8278_cse , and_8286_cse , and_8295_cse , and_8305_cse , and_8316_cse
          , and_8328_cse , and_8341_cse , and_8355_cse , and_8362_cse});
      reg_div_mgc_div_8_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_65_sg1
          , delta_conc_3_tmp_mut_66_sg1 , delta_conc_3_tmp_mut_67_sg1 , delta_conc_3_tmp_mut_68_sg1
          , delta_conc_3_tmp_mut_69_sg1 , delta_conc_3_tmp_mut_70_sg1 , delta_conc_3_tmp_mut_71_sg1
          , delta_conc_3_tmp_mut_72_sg1}, {and_8457_cse , and_8465_cse , and_8474_cse
          , and_8484_cse , and_8495_cse , and_8507_cse , and_8520_cse , and_8534_cse
          , and_8541_cse});
      reg_div_mgc_div_8_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_65_sg1 , else_7_else_1_else_conc_tmp_mut_66_sg1
          , else_7_else_1_else_conc_tmp_mut_67_sg1 , else_7_else_1_else_conc_tmp_mut_68_sg1
          , else_7_else_1_else_conc_tmp_mut_69_sg1 , else_7_else_1_else_conc_tmp_mut_70_sg1
          , else_7_else_1_else_conc_tmp_mut_71_sg1 , else_7_else_1_else_conc_tmp_mut_72_sg1},
          {and_8457_cse , and_8465_cse , and_8474_cse , and_8484_cse , and_8495_cse
          , and_8507_cse , and_8520_cse , and_8534_cse , and_8541_cse});
      reg_div_mgc_div_9_b_tmp <= MUX1HOT_v_16_9_2({(else_7_acc_3_itm[16:1]) , delta_conc_3_tmp_mut_73_sg1
          , delta_conc_3_tmp_mut_74_sg1 , delta_conc_3_tmp_mut_75_sg1 , delta_conc_3_tmp_mut_76_sg1
          , delta_conc_3_tmp_mut_77_sg1 , delta_conc_3_tmp_mut_78_sg1 , delta_conc_3_tmp_mut_79_sg1
          , delta_conc_3_tmp_mut_80_sg1}, {and_8636_cse , and_8644_cse , and_8653_cse
          , and_8663_cse , and_8673_cse , and_8682_cse , and_8691_cse , and_8700_cse
          , and_8702_cse});
      reg_div_mgc_div_9_a_tmp <= MUX1HOT_v_17_9_2({(else_7_else_1_else_acc_2_itm[17:1])
          , else_7_else_1_else_conc_tmp_mut_73_sg1 , else_7_else_1_else_conc_tmp_mut_74_sg1
          , else_7_else_1_else_conc_tmp_mut_75_sg1 , else_7_else_1_else_conc_tmp_mut_76_sg1
          , else_7_else_1_else_conc_tmp_mut_77_sg1 , else_7_else_1_else_conc_tmp_mut_78_sg1
          , else_7_else_1_else_conc_tmp_mut_79_sg1 , else_7_else_1_else_conc_tmp_mut_80_sg1},
          {and_8636_cse , and_8644_cse , and_8653_cse , and_8663_cse , and_8673_cse
          , and_8682_cse , and_8691_cse , and_8700_cse , and_8702_cse});
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [1:0] inputs;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[1:1];
      end
      1'b1 : begin
        result = inputs[0:0];
      end
      default : begin
        result = inputs[1:1];
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [15:0] MUX_v_16_2_2;
    input [31:0] inputs;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[31:16];
      end
      1'b1 : begin
        result = inputs[15:0];
      end
      default : begin
        result = inputs[31:16];
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function [29:0] MUX1HOT_v_30_10_2;
    input [299:0] inputs;
    input [9:0] sel;
    reg [29:0] result;
    integer i;
  begin
    result = inputs[0+:30] & {30{sel[0]}};
    for( i = 1; i < 10; i = i + 1 )
      result = result | (inputs[i*30+:30] & {30{sel[i]}});
    MUX1HOT_v_30_10_2 = result;
  end
  endfunction


  function [12:0] MUX1HOT_v_13_10_2;
    input [129:0] inputs;
    input [9:0] sel;
    reg [12:0] result;
    integer i;
  begin
    result = inputs[0+:13] & {13{sel[0]}};
    for( i = 1; i < 10; i = i + 1 )
      result = result | (inputs[i*13+:13] & {13{sel[i]}});
    MUX1HOT_v_13_10_2 = result;
  end
  endfunction


  function [11:0] MUX1HOT_v_12_3_2;
    input [35:0] inputs;
    input [2:0] sel;
    reg [11:0] result;
    integer i;
  begin
    result = inputs[0+:12] & {12{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*12+:12] & {12{sel[i]}});
    MUX1HOT_v_12_3_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [2:0] inputs;
    input [2:0] sel;
    reg [0:0] result;
    integer i;
  begin
    result = inputs[0+:1] & {1{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*1+:1] & {1{sel[i]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [16:0] MUX1HOT_v_17_12_2;
    input [203:0] inputs;
    input [11:0] sel;
    reg [16:0] result;
    integer i;
  begin
    result = inputs[0+:17] & {17{sel[0]}};
    for( i = 1; i < 12; i = i + 1 )
      result = result | (inputs[i*17+:17] & {17{sel[i]}});
    MUX1HOT_v_17_12_2 = result;
  end
  endfunction


  function [15:0] MUX1HOT_v_16_3_2;
    input [47:0] inputs;
    input [2:0] sel;
    reg [15:0] result;
    integer i;
  begin
    result = inputs[0+:16] & {16{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*16+:16] & {16{sel[i]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [63:0] inputs;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[63:32];
      end
      1'b1 : begin
        result = inputs[31:0];
      end
      default : begin
        result = inputs[63:32];
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [15:0] MUX1HOT_v_16_10_2;
    input [159:0] inputs;
    input [9:0] sel;
    reg [15:0] result;
    integer i;
  begin
    result = inputs[0+:16] & {16{sel[0]}};
    for( i = 1; i < 10; i = i + 1 )
      result = result | (inputs[i*16+:16] & {16{sel[i]}});
    MUX1HOT_v_16_10_2 = result;
  end
  endfunction


  function [15:0] signext_16_1;
    input [0:0] vector;
  begin
    signext_16_1= {{15{vector[0]}}, vector};
  end
  endfunction


  function [29:0] signext_30_21;
    input [20:0] vector;
  begin
    signext_30_21= {{9{vector[20]}}, vector};
  end
  endfunction


  function [12:0] MUX_v_13_2_2;
    input [25:0] inputs;
    input [0:0] sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[25:13];
      end
      1'b1 : begin
        result = inputs[12:0];
      end
      default : begin
        result = inputs[25:13];
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function [12:0] signext_13_1;
    input [0:0] vector;
  begin
    signext_13_1= {{12{vector[0]}}, vector};
  end
  endfunction


  function [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function [31:0] signext_32_16;
    input [15:0] vector;
  begin
    signext_32_16= {{16{vector[15]}}, vector};
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [7:0] inputs;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[7:4];
      end
      1'b1 : begin
        result = inputs[3:0];
      end
      default : begin
        result = inputs[7:4];
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [16:0] MUX_v_17_2_2;
    input [33:0] inputs;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[33:17];
      end
      1'b1 : begin
        result = inputs[16:0];
      end
      default : begin
        result = inputs[33:17];
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function [14:0] readslicef_69_15_54;
    input [68:0] vector;
    reg [68:0] tmp;
  begin
    tmp = vector >> 54;
    readslicef_69_15_54 = tmp[14:0];
  end
  endfunction


  function [15:0] MUX1HOT_v_16_9_2;
    input [143:0] inputs;
    input [8:0] sel;
    reg [15:0] result;
    integer i;
  begin
    result = inputs[0+:16] & {16{sel[0]}};
    for( i = 1; i < 9; i = i + 1 )
      result = result | (inputs[i*16+:16] & {16{sel[i]}});
    MUX1HOT_v_16_9_2 = result;
  end
  endfunction


  function [16:0] MUX1HOT_v_17_9_2;
    input [152:0] inputs;
    input [8:0] sel;
    reg [16:0] result;
    integer i;
  begin
    result = inputs[0+:17] & {17{sel[0]}};
    for( i = 1; i < 9; i = i + 1 )
      result = result | (inputs[i*17+:17] & {17{sel[i]}});
    MUX1HOT_v_17_9_2 = result;
  end
  endfunction


  function  [17:0] conv_s2u_17_18 ;
    input signed [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function  [3:0] conv_u2u_1_4 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_4 = {{3{1'b0}}, vector};
  end
  endfunction


  function  [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function signed [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 = {1'b0, vector};
  end
  endfunction


  function  [20:0] conv_s2u_42_21 ;
    input signed [41:0]  vector ;
  begin
    conv_s2u_42_21 = vector[20:0];
  end
  endfunction


  function signed [20:0] conv_s2s_16_21 ;
    input signed [15:0]  vector ;
  begin
    conv_s2s_16_21 = {{5{vector[15]}}, vector};
  end
  endfunction


  function  [68:0] conv_s2u_138_69 ;
    input signed [137:0]  vector ;
  begin
    conv_s2u_138_69 = vector[68:0];
  end
  endfunction


  function signed [68:0] conv_s2s_16_69 ;
    input signed [15:0]  vector ;
  begin
    conv_s2s_16_69 = {{53{vector[15]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HSVRGB
//  Generated from file(s):
//    2) $PROJECT_HOME/../RGBHSV/RGBHSV.cpp
// ------------------------------------------------------------------


module HSVRGB (
  R_IN_rsc_z, G_IN_rsc_z, B_IN_rsc_z, H_OUT_rsc_z, S_OUT_rsc_z, V_OUT_rsc_z, clk,
      rst
);
  input [31:0] R_IN_rsc_z;
  input [31:0] G_IN_rsc_z;
  input [31:0] B_IN_rsc_z;
  output [31:0] H_OUT_rsc_z;
  output [31:0] S_OUT_rsc_z;
  output [31:0] V_OUT_rsc_z;
  input clk;
  input rst;


  // Interconnect Declarations
  wire [31:0] R_IN_rsc_mgc_in_wire_d;
  wire [31:0] G_IN_rsc_mgc_in_wire_d;
  wire [31:0] B_IN_rsc_mgc_in_wire_d;
  wire [31:0] H_OUT_rsc_mgc_out_stdreg_d;
  wire [31:0] S_OUT_rsc_mgc_out_stdreg_d;
  wire [31:0] V_OUT_rsc_mgc_out_stdreg_d;
  wire [48:0] div_mgc_div_a;
  wire [31:0] div_mgc_div_b;
  wire [48:0] div_mgc_div_z;
  wire [48:0] div_mgc_div_1_a;
  wire [31:0] div_mgc_div_1_b;
  wire [48:0] div_mgc_div_1_z;
  wire [48:0] div_mgc_div_2_a;
  wire [31:0] div_mgc_div_2_b;
  wire [48:0] div_mgc_div_2_z;
  wire [48:0] div_mgc_div_3_a;
  wire [31:0] div_mgc_div_3_b;
  wire [48:0] div_mgc_div_3_z;
  wire [48:0] div_mgc_div_4_a;
  wire [31:0] div_mgc_div_4_b;
  wire [48:0] div_mgc_div_4_z;
  wire [48:0] div_mgc_div_5_a;
  wire [31:0] div_mgc_div_5_b;
  wire [48:0] div_mgc_div_5_z;
  wire [48:0] div_mgc_div_6_a;
  wire [31:0] div_mgc_div_6_b;
  wire [48:0] div_mgc_div_6_z;
  wire [48:0] div_mgc_div_7_a;
  wire [31:0] div_mgc_div_7_b;
  wire [48:0] div_mgc_div_7_z;
  wire [48:0] div_mgc_div_8_a;
  wire [31:0] div_mgc_div_8_b;
  wire [48:0] div_mgc_div_8_z;
  wire [48:0] div_mgc_div_9_a;
  wire [31:0] div_mgc_div_9_b;
  wire [48:0] div_mgc_div_9_z;
  wire [48:0] div_mgc_div_10_a;
  wire [31:0] div_mgc_div_10_b;
  wire [48:0] div_mgc_div_10_z;
  wire [48:0] div_mgc_div_11_a;
  wire [31:0] div_mgc_div_11_b;
  wire [48:0] div_mgc_div_11_z;
  wire [48:0] div_mgc_div_12_a;
  wire [31:0] div_mgc_div_12_b;
  wire [48:0] div_mgc_div_12_z;
  wire [48:0] div_mgc_div_13_a;
  wire [31:0] div_mgc_div_13_b;
  wire [48:0] div_mgc_div_13_z;
  wire [48:0] div_mgc_div_14_a;
  wire [31:0] div_mgc_div_14_b;
  wire [48:0] div_mgc_div_14_z;
  wire [48:0] div_mgc_div_15_a;
  wire [31:0] div_mgc_div_15_b;
  wire [48:0] div_mgc_div_15_z;
  wire [48:0] div_mgc_div_16_a;
  wire [31:0] div_mgc_div_16_b;
  wire [48:0] div_mgc_div_16_z;
  wire [48:0] div_mgc_div_17_a;
  wire [31:0] div_mgc_div_17_b;
  wire [48:0] div_mgc_div_17_z;
  wire [48:0] div_mgc_div_18_a;
  wire [31:0] div_mgc_div_18_b;
  wire [48:0] div_mgc_div_18_z;
  wire [48:0] div_mgc_div_19_a;
  wire [31:0] div_mgc_div_19_b;
  wire [48:0] div_mgc_div_19_z;
  wire [48:0] div_mgc_div_20_a;
  wire [31:0] div_mgc_div_20_b;
  wire [48:0] div_mgc_div_20_z;
  wire [48:0] div_mgc_div_21_a;
  wire [31:0] div_mgc_div_21_b;
  wire [48:0] div_mgc_div_21_z;
  wire [48:0] div_mgc_div_22_a;
  wire [31:0] div_mgc_div_22_b;
  wire [48:0] div_mgc_div_22_z;
  wire [48:0] div_mgc_div_23_a;
  wire [31:0] div_mgc_div_23_b;
  wire [48:0] div_mgc_div_23_z;
  wire [48:0] div_mgc_div_24_a;
  wire [31:0] div_mgc_div_24_b;
  wire [48:0] div_mgc_div_24_z;
  wire [48:0] div_mgc_div_25_a;
  wire [31:0] div_mgc_div_25_b;
  wire [48:0] div_mgc_div_25_z;
  wire [48:0] div_mgc_div_26_a;
  wire [31:0] div_mgc_div_26_b;
  wire [48:0] div_mgc_div_26_z;
  wire [47:0] div_mgc_div_27_a;
  wire [31:0] div_mgc_div_27_b;
  wire [47:0] div_mgc_div_27_z;
  wire [47:0] div_mgc_div_28_a;
  wire [31:0] div_mgc_div_28_b;
  wire [47:0] div_mgc_div_28_z;
  wire [47:0] div_mgc_div_29_a;
  wire [31:0] div_mgc_div_29_b;
  wire [47:0] div_mgc_div_29_z;
  wire [47:0] div_mgc_div_30_a;
  wire [31:0] div_mgc_div_30_b;
  wire [47:0] div_mgc_div_30_z;
  wire [47:0] div_mgc_div_31_a;
  wire [31:0] div_mgc_div_31_b;
  wire [47:0] div_mgc_div_31_z;
  wire [47:0] div_mgc_div_32_a;
  wire [31:0] div_mgc_div_32_b;
  wire [47:0] div_mgc_div_32_z;
  wire [47:0] div_mgc_div_33_a;
  wire [31:0] div_mgc_div_33_b;
  wire [47:0] div_mgc_div_33_z;
  wire [47:0] div_mgc_div_34_a;
  wire [31:0] div_mgc_div_34_b;
  wire [47:0] div_mgc_div_34_z;
  wire [47:0] div_mgc_div_35_a;
  wire [31:0] div_mgc_div_35_b;
  wire [47:0] div_mgc_div_35_z;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire #(.rscid(1),
  .width(32)) R_IN_rsc_mgc_in_wire (
      .d(R_IN_rsc_mgc_in_wire_d),
      .z(R_IN_rsc_z)
    );
  mgc_in_wire #(.rscid(2),
  .width(32)) G_IN_rsc_mgc_in_wire (
      .d(G_IN_rsc_mgc_in_wire_d),
      .z(G_IN_rsc_z)
    );
  mgc_in_wire #(.rscid(3),
  .width(32)) B_IN_rsc_mgc_in_wire (
      .d(B_IN_rsc_mgc_in_wire_d),
      .z(B_IN_rsc_z)
    );
  mgc_out_stdreg #(.rscid(4),
  .width(32)) H_OUT_rsc_mgc_out_stdreg (
      .d(H_OUT_rsc_mgc_out_stdreg_d),
      .z(H_OUT_rsc_z)
    );
  mgc_out_stdreg #(.rscid(5),
  .width(32)) S_OUT_rsc_mgc_out_stdreg (
      .d(S_OUT_rsc_mgc_out_stdreg_d),
      .z(S_OUT_rsc_z)
    );
  mgc_out_stdreg #(.rscid(6),
  .width(32)) V_OUT_rsc_mgc_out_stdreg (
      .d(V_OUT_rsc_mgc_out_stdreg_d),
      .z(V_OUT_rsc_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div (
      .a(div_mgc_div_a),
      .b(div_mgc_div_b),
      .z(div_mgc_div_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_1 (
      .a(div_mgc_div_1_a),
      .b(div_mgc_div_1_b),
      .z(div_mgc_div_1_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_2 (
      .a(div_mgc_div_2_a),
      .b(div_mgc_div_2_b),
      .z(div_mgc_div_2_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_3 (
      .a(div_mgc_div_3_a),
      .b(div_mgc_div_3_b),
      .z(div_mgc_div_3_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_4 (
      .a(div_mgc_div_4_a),
      .b(div_mgc_div_4_b),
      .z(div_mgc_div_4_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_5 (
      .a(div_mgc_div_5_a),
      .b(div_mgc_div_5_b),
      .z(div_mgc_div_5_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_6 (
      .a(div_mgc_div_6_a),
      .b(div_mgc_div_6_b),
      .z(div_mgc_div_6_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_7 (
      .a(div_mgc_div_7_a),
      .b(div_mgc_div_7_b),
      .z(div_mgc_div_7_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_8 (
      .a(div_mgc_div_8_a),
      .b(div_mgc_div_8_b),
      .z(div_mgc_div_8_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_9 (
      .a(div_mgc_div_9_a),
      .b(div_mgc_div_9_b),
      .z(div_mgc_div_9_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_10 (
      .a(div_mgc_div_10_a),
      .b(div_mgc_div_10_b),
      .z(div_mgc_div_10_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_11 (
      .a(div_mgc_div_11_a),
      .b(div_mgc_div_11_b),
      .z(div_mgc_div_11_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_12 (
      .a(div_mgc_div_12_a),
      .b(div_mgc_div_12_b),
      .z(div_mgc_div_12_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_13 (
      .a(div_mgc_div_13_a),
      .b(div_mgc_div_13_b),
      .z(div_mgc_div_13_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_14 (
      .a(div_mgc_div_14_a),
      .b(div_mgc_div_14_b),
      .z(div_mgc_div_14_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_15 (
      .a(div_mgc_div_15_a),
      .b(div_mgc_div_15_b),
      .z(div_mgc_div_15_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_16 (
      .a(div_mgc_div_16_a),
      .b(div_mgc_div_16_b),
      .z(div_mgc_div_16_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_17 (
      .a(div_mgc_div_17_a),
      .b(div_mgc_div_17_b),
      .z(div_mgc_div_17_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_18 (
      .a(div_mgc_div_18_a),
      .b(div_mgc_div_18_b),
      .z(div_mgc_div_18_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_19 (
      .a(div_mgc_div_19_a),
      .b(div_mgc_div_19_b),
      .z(div_mgc_div_19_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_20 (
      .a(div_mgc_div_20_a),
      .b(div_mgc_div_20_b),
      .z(div_mgc_div_20_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_21 (
      .a(div_mgc_div_21_a),
      .b(div_mgc_div_21_b),
      .z(div_mgc_div_21_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_22 (
      .a(div_mgc_div_22_a),
      .b(div_mgc_div_22_b),
      .z(div_mgc_div_22_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_23 (
      .a(div_mgc_div_23_a),
      .b(div_mgc_div_23_b),
      .z(div_mgc_div_23_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_24 (
      .a(div_mgc_div_24_a),
      .b(div_mgc_div_24_b),
      .z(div_mgc_div_24_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_25 (
      .a(div_mgc_div_25_a),
      .b(div_mgc_div_25_b),
      .z(div_mgc_div_25_z)
    );
  mgc_div #(.width_a(49),
  .width_b(32),
  .signd(1)) div_mgc_div_26 (
      .a(div_mgc_div_26_a),
      .b(div_mgc_div_26_b),
      .z(div_mgc_div_26_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_27 (
      .a(div_mgc_div_27_a),
      .b(div_mgc_div_27_b),
      .z(div_mgc_div_27_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_28 (
      .a(div_mgc_div_28_a),
      .b(div_mgc_div_28_b),
      .z(div_mgc_div_28_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_29 (
      .a(div_mgc_div_29_a),
      .b(div_mgc_div_29_b),
      .z(div_mgc_div_29_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_30 (
      .a(div_mgc_div_30_a),
      .b(div_mgc_div_30_b),
      .z(div_mgc_div_30_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_31 (
      .a(div_mgc_div_31_a),
      .b(div_mgc_div_31_b),
      .z(div_mgc_div_31_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_32 (
      .a(div_mgc_div_32_a),
      .b(div_mgc_div_32_b),
      .z(div_mgc_div_32_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_33 (
      .a(div_mgc_div_33_a),
      .b(div_mgc_div_33_b),
      .z(div_mgc_div_33_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_34 (
      .a(div_mgc_div_34_a),
      .b(div_mgc_div_34_b),
      .z(div_mgc_div_34_z)
    );
  mgc_div #(.width_a(48),
  .width_b(32),
  .signd(1)) div_mgc_div_35 (
      .a(div_mgc_div_35_a),
      .b(div_mgc_div_35_b),
      .z(div_mgc_div_35_z)
    );
  HSVRGB_core HSVRGB_core_inst (
      .clk(clk),
      .rst(rst),
      .R_IN_rsc_mgc_in_wire_d(R_IN_rsc_mgc_in_wire_d),
      .G_IN_rsc_mgc_in_wire_d(G_IN_rsc_mgc_in_wire_d),
      .B_IN_rsc_mgc_in_wire_d(B_IN_rsc_mgc_in_wire_d),
      .H_OUT_rsc_mgc_out_stdreg_d(H_OUT_rsc_mgc_out_stdreg_d),
      .S_OUT_rsc_mgc_out_stdreg_d(S_OUT_rsc_mgc_out_stdreg_d),
      .V_OUT_rsc_mgc_out_stdreg_d(V_OUT_rsc_mgc_out_stdreg_d),
      .div_mgc_div_a(div_mgc_div_a),
      .div_mgc_div_b(div_mgc_div_b),
      .div_mgc_div_z(div_mgc_div_z),
      .div_mgc_div_1_a(div_mgc_div_1_a),
      .div_mgc_div_1_b(div_mgc_div_1_b),
      .div_mgc_div_1_z(div_mgc_div_1_z),
      .div_mgc_div_2_a(div_mgc_div_2_a),
      .div_mgc_div_2_b(div_mgc_div_2_b),
      .div_mgc_div_2_z(div_mgc_div_2_z),
      .div_mgc_div_3_a(div_mgc_div_3_a),
      .div_mgc_div_3_b(div_mgc_div_3_b),
      .div_mgc_div_3_z(div_mgc_div_3_z),
      .div_mgc_div_4_a(div_mgc_div_4_a),
      .div_mgc_div_4_b(div_mgc_div_4_b),
      .div_mgc_div_4_z(div_mgc_div_4_z),
      .div_mgc_div_5_a(div_mgc_div_5_a),
      .div_mgc_div_5_b(div_mgc_div_5_b),
      .div_mgc_div_5_z(div_mgc_div_5_z),
      .div_mgc_div_6_a(div_mgc_div_6_a),
      .div_mgc_div_6_b(div_mgc_div_6_b),
      .div_mgc_div_6_z(div_mgc_div_6_z),
      .div_mgc_div_7_a(div_mgc_div_7_a),
      .div_mgc_div_7_b(div_mgc_div_7_b),
      .div_mgc_div_7_z(div_mgc_div_7_z),
      .div_mgc_div_8_a(div_mgc_div_8_a),
      .div_mgc_div_8_b(div_mgc_div_8_b),
      .div_mgc_div_8_z(div_mgc_div_8_z),
      .div_mgc_div_9_a(div_mgc_div_9_a),
      .div_mgc_div_9_b(div_mgc_div_9_b),
      .div_mgc_div_9_z(div_mgc_div_9_z),
      .div_mgc_div_10_a(div_mgc_div_10_a),
      .div_mgc_div_10_b(div_mgc_div_10_b),
      .div_mgc_div_10_z(div_mgc_div_10_z),
      .div_mgc_div_11_a(div_mgc_div_11_a),
      .div_mgc_div_11_b(div_mgc_div_11_b),
      .div_mgc_div_11_z(div_mgc_div_11_z),
      .div_mgc_div_12_a(div_mgc_div_12_a),
      .div_mgc_div_12_b(div_mgc_div_12_b),
      .div_mgc_div_12_z(div_mgc_div_12_z),
      .div_mgc_div_13_a(div_mgc_div_13_a),
      .div_mgc_div_13_b(div_mgc_div_13_b),
      .div_mgc_div_13_z(div_mgc_div_13_z),
      .div_mgc_div_14_a(div_mgc_div_14_a),
      .div_mgc_div_14_b(div_mgc_div_14_b),
      .div_mgc_div_14_z(div_mgc_div_14_z),
      .div_mgc_div_15_a(div_mgc_div_15_a),
      .div_mgc_div_15_b(div_mgc_div_15_b),
      .div_mgc_div_15_z(div_mgc_div_15_z),
      .div_mgc_div_16_a(div_mgc_div_16_a),
      .div_mgc_div_16_b(div_mgc_div_16_b),
      .div_mgc_div_16_z(div_mgc_div_16_z),
      .div_mgc_div_17_a(div_mgc_div_17_a),
      .div_mgc_div_17_b(div_mgc_div_17_b),
      .div_mgc_div_17_z(div_mgc_div_17_z),
      .div_mgc_div_18_a(div_mgc_div_18_a),
      .div_mgc_div_18_b(div_mgc_div_18_b),
      .div_mgc_div_18_z(div_mgc_div_18_z),
      .div_mgc_div_19_a(div_mgc_div_19_a),
      .div_mgc_div_19_b(div_mgc_div_19_b),
      .div_mgc_div_19_z(div_mgc_div_19_z),
      .div_mgc_div_20_a(div_mgc_div_20_a),
      .div_mgc_div_20_b(div_mgc_div_20_b),
      .div_mgc_div_20_z(div_mgc_div_20_z),
      .div_mgc_div_21_a(div_mgc_div_21_a),
      .div_mgc_div_21_b(div_mgc_div_21_b),
      .div_mgc_div_21_z(div_mgc_div_21_z),
      .div_mgc_div_22_a(div_mgc_div_22_a),
      .div_mgc_div_22_b(div_mgc_div_22_b),
      .div_mgc_div_22_z(div_mgc_div_22_z),
      .div_mgc_div_23_a(div_mgc_div_23_a),
      .div_mgc_div_23_b(div_mgc_div_23_b),
      .div_mgc_div_23_z(div_mgc_div_23_z),
      .div_mgc_div_24_a(div_mgc_div_24_a),
      .div_mgc_div_24_b(div_mgc_div_24_b),
      .div_mgc_div_24_z(div_mgc_div_24_z),
      .div_mgc_div_25_a(div_mgc_div_25_a),
      .div_mgc_div_25_b(div_mgc_div_25_b),
      .div_mgc_div_25_z(div_mgc_div_25_z),
      .div_mgc_div_26_a(div_mgc_div_26_a),
      .div_mgc_div_26_b(div_mgc_div_26_b),
      .div_mgc_div_26_z(div_mgc_div_26_z),
      .div_mgc_div_27_a(div_mgc_div_27_a),
      .div_mgc_div_27_b(div_mgc_div_27_b),
      .div_mgc_div_27_z(div_mgc_div_27_z),
      .div_mgc_div_28_a(div_mgc_div_28_a),
      .div_mgc_div_28_b(div_mgc_div_28_b),
      .div_mgc_div_28_z(div_mgc_div_28_z),
      .div_mgc_div_29_a(div_mgc_div_29_a),
      .div_mgc_div_29_b(div_mgc_div_29_b),
      .div_mgc_div_29_z(div_mgc_div_29_z),
      .div_mgc_div_30_a(div_mgc_div_30_a),
      .div_mgc_div_30_b(div_mgc_div_30_b),
      .div_mgc_div_30_z(div_mgc_div_30_z),
      .div_mgc_div_31_a(div_mgc_div_31_a),
      .div_mgc_div_31_b(div_mgc_div_31_b),
      .div_mgc_div_31_z(div_mgc_div_31_z),
      .div_mgc_div_32_a(div_mgc_div_32_a),
      .div_mgc_div_32_b(div_mgc_div_32_b),
      .div_mgc_div_32_z(div_mgc_div_32_z),
      .div_mgc_div_33_a(div_mgc_div_33_a),
      .div_mgc_div_33_b(div_mgc_div_33_b),
      .div_mgc_div_33_z(div_mgc_div_33_z),
      .div_mgc_div_34_a(div_mgc_div_34_a),
      .div_mgc_div_34_b(div_mgc_div_34_b),
      .div_mgc_div_34_z(div_mgc_div_34_z),
      .div_mgc_div_35_a(div_mgc_div_35_a),
      .div_mgc_div_35_b(div_mgc_div_35_b),
      .div_mgc_div_35_z(div_mgc_div_35_z)
    );
endmodule



