library verilog;
use verilog.vl_types.all;
entity MazeRAMTester_vlg_vec_tst is
end MazeRAMTester_vlg_vec_tst;
