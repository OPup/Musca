library verilog;
use verilog.vl_types.all;
entity MazeRAMTester_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end MazeRAMTester_vlg_sample_tst;
