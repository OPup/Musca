
//------> ./rtl_mgc_ioport.v 
//------------------------------------------------------------------
//                M G C _ I O P O R T _ C O M P S
//------------------------------------------------------------------

//------------------------------------------------------------------
//                       M O D U L E S
//------------------------------------------------------------------

//------------------------------------------------------------------
//-- INPUT ENTITIES
//------------------------------------------------------------------

module mgc_in_wire (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output [width-1:0] d;
  output             lz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule
//------------------------------------------------------------------

module mgc_chan_in (ld, vd, d, lz, vz, z, size, req_size, sizez, sizelz);

  parameter integer rscid = 1;
  parameter integer width = 8;
  parameter integer sz_width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;
  output [sz_width-1:0] size;
  input              req_size;
  input  [sz_width-1:0] sizez;
  output             sizelz;


  wire               vd;
  wire   [width-1:0] d;
  wire               lz;
  wire   [sz_width-1:0] size;
  wire               sizelz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;
  assign size = sizez;
  assign sizelz = req_size;

endmodule


//------------------------------------------------------------------
//-- OUTPUT ENTITIES
//------------------------------------------------------------------

module mgc_out_stdreg (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  input  [width-1:0] d;
  output             lz;
  output [width-1:0] z;

  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_out_prereg_en (ld, d, lz, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    wire               lz;
    wire   [width-1:0] z;

    assign z = d;
    assign lz = ld;

endmodule

//------------------------------------------------------------------
//-- INOUT ENTITIES
//------------------------------------------------------------------

module mgc_inout_stdreg_en (ldin, din, ldout, dout, lzin, lzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    output             lzin;
    output             lzout;
    inout  [width-1:0] z;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign z = ldout ? dout : {width{1'bz}};

endmodule

//------------------------------------------------------------------
module hid_tribuf( I_SIG, ENABLE, O_SIG);
  parameter integer width = 8;

  input [width-1:0] I_SIG;
  input ENABLE;
  inout [width-1:0] O_SIG;

  assign O_SIG = (ENABLE) ? I_SIG : { width{1'bz}};

endmodule
//------------------------------------------------------------------

module mgc_inout_stdreg_wait (ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;
    wire   ldout_and_vzout;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign vdout = vzout ;
    assign ldout_and_vzout = ldout && vzout ;

    hid_tribuf #(width) tb( .I_SIG(dout),
                            .ENABLE(ldout_and_vzout),
                            .O_SIG(z) );

endmodule

//------------------------------------------------------------------

module mgc_inout_buf_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    hid_tribuf #(width) tb( .I_SIG(z_buf),
                            .ENABLE((lzout_buf && (!ldin) && vzout) ),
                            .O_SIG(z)  );

    mgc_out_buf_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFF
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );


endmodule

module mgc_inout_fifo_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer ph_log2 = 3;     // log2(fifo_sz)
    parameter integer pwropt  = 0;     // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               comb;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    assign comb = (lzout_buf && (!ldin) && vzout);

    hid_tribuf #(width) tb2( .I_SIG(z_buf), .ENABLE(comb), .O_SIG(z)  );

    mgc_out_fifo_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
    )
    FIFO
    (
        .clk   (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );

endmodule

//------------------------------------------------------------------
//-- I/O SYNCHRONIZATION ENTITIES
//------------------------------------------------------------------

module mgc_io_sync (ld, lz);

    input  ld;
    output lz;

    assign lz = ld;

endmodule

module mgc_bsync_rdy (rd, rz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 0;

    input  rd;
    output rz;

    wire   rz;

    assign rz = rd;

endmodule

module mgc_bsync_vld (vd, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 0;
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule

module mgc_bsync_rv (rd, vd, rz, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 1;

    input  rd;
    output vd;
    output rz;
    input  vz;

    wire   vd;
    wire   rz;

    assign rz = rd;
    assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_sync (ldin, vdin, ldout, vdout);

  input  ldin;
  output vdin;
  input  ldout;
  output vdout;

  wire   vdin;
  wire   vdout;

  assign vdin = ldout;
  assign vdout = ldin;

endmodule

///////////////////////////////////////////////////////////////////////////////
// dummy function used to preserve funccalls for modulario
// it looks like a memory read to the caller
///////////////////////////////////////////////////////////////////////////////
module funccall_inout (d, ad, bd, z, az, bz);

  parameter integer ram_id = 1;
  parameter integer width = 8;
  parameter integer addr_width = 8;

  output [width-1:0]       d;
  input  [addr_width-1:0]  ad;
  input                    bd;
  input  [width-1:0]       z;
  output [addr_width-1:0]  az;
  output                   bz;

  wire   [width-1:0]       d;
  wire   [addr_width-1:0]  az;
  wire                     bz;

  assign d  = z;
  assign az = ad;
  assign bz = bd;

endmodule


///////////////////////////////////////////////////////////////////////////////
// inlinable modular io not otherwise found in mgc_ioport
///////////////////////////////////////////////////////////////////////////////

module modulario_en_in (vd, d, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output             vd;
  output [width-1:0] d;
  input              vz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               vd;

  assign d = z;
  assign vd = vz;

endmodule

//------> ./rtl_mgc_ioport_v2001.v 
//------------------------------------------------------------------

module mgc_out_reg_pos (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(posedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(posedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg_neg (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(negedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(negedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg (clk, en, arst, srst, ld, d, lz, z); // Not Supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;


    generate
    if (ph_clk == 1'b0)
    begin: NEG_EDGE

        mgc_out_reg_neg
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_neg_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    else
    begin: POS_EDGE

        mgc_out_reg_pos
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_pos_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    endgenerate

endmodule




//------------------------------------------------------------------

module mgc_out_buf_wait (clk, en, arst, srst, ld, vd, d, vz, lz, z); // Not supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    output             vd;
    input  [width-1:0] d;
    output             lz;
    input              vz;
    output [width-1:0] z;

    wire               filled;
    wire               filled_next;
    wire   [width-1:0] abuf;
    wire               lbuf;


    assign filled_next = (filled & (~vz)) | (filled & ld) | (ld & (~vz));

    assign lbuf = ld & ~(filled ^ vz);

    assign vd = vz | ~filled;

    assign lz = ld | filled;

    assign z = (filled) ? abuf : d;

    wire dummy;
    wire dummy_bufreg_lz;

    // Output registers:
    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (1'b1),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    STATREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (filled_next),
        .d       (1'b0),       // input d is unused
        .lz      (filled),
        .z       (dummy)            // output z is unused
    );

    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (lbuf),
        .d       (d),
        .lz      (dummy_bufreg_lz),
        .z       (abuf)
    );

endmodule

//------------------------------------------------------------------

module mgc_out_fifo_wait (clk, en, arst, srst, ld, vd, d, lz, vz,  z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1; // clock enable polarity
    parameter         ph_arst = 1'b1; // async reset polarity
    parameter         ph_srst = 1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt


    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;

    wire    [31:0]      size;


      // Output registers:
 mgc_out_fifo_wait_core#(
        .rscid   (rscid),
        .width   (width),
        .sz_width (32),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
        ) CORE (
        .clk (clk),
        .en (en),
        .arst (arst),
        .srst (srst),
        .ld (ld),
        .vd (vd),
        .d (d),
        .lz (lz),
        .vz (vz),
        .z (z),
        .size (size)
        );

endmodule



module mgc_out_fifo_wait_core (clk, en, arst, srst, ld, vd, d, lz, vz,  z, size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // size of port for elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt

   localparam integer  fifo_b = width * fifo_sz;

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;
    output    [sz_width-1:0]      size;

    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat_pre;
    wire     [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] en_l;
    reg      [(((fifo_sz > 0) ? fifo_sz : 1)-1)/8:0] en_l_s;

    reg       [width-1:0] buff_nxt;

    reg                   stat_nxt;
    reg                   stat_before;
    reg                   stat_after;
    reg                   en_l_var;

    integer               i;
    genvar                eni;

    wire [32:0]           size_t;
    reg [31:0]            count;
    reg [31:0]            count_t;
    reg [32:0]            n_elem;
// pragma translate_off
    reg [31:0]            peak;
// pragma translate_on

    wire [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] dummy_statreg_lz;
    wire [( (fifo_b > 0) ? fifo_b : 1)-1:0] dummy_bufreg_lz;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      assign vd = vz | ~stat[0];
      assign lz = ld | stat[fifo_sz-1];
      assign size_t = (count - (vz && stat[fifo_sz-1])) + ld;
      assign size = size_t[sz_width-1:0];
      assign z = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : d;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          if (i != 0)
            stat_before = stat[i-1];
          else
            stat_before = 1'b0;

          if (i != (fifo_sz-1))
            stat_after = stat[i+1];
          else
            stat_after = 1'b1;

          stat_nxt = stat_after &
                    (stat_before | (stat[i] & (~vz)) | (stat[i] & ld) | (ld & (~vz)));

          stat_pre[i] = stat_nxt;
          en_l_var = 1'b1;
          if (!stat_nxt)
            begin
              buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end
          else if (vz && stat_before)
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
          else if (ld && !((vz && stat_before) || ((!vz) && stat[i])))
            buff_nxt = d;
          else
            begin
              if (pwropt == 0)
                buff_nxt[0+:width] = buff[width*i+:width];
              else
                buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if ((stat_after == 1'b1) && (stat[i] == 1'b0))
            n_elem = ($unsigned(fifo_sz) - 1) - i;
        end

        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b1;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b0;

        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if ((i%'d2) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]|stat_pre[i-1]);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]|stat_pre[i-1]);
          end
        end

        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = { {(32-ph_log2){1'b0}}, fifo_sz};
        else
          count_t = n_elem[31:0];
        count = count_t;
// pragma translate_off
        if ( peak < count )
          peak = count;
// pragma translate_on
      end

      if (pwropt == 0)
      begin: NOCGFIFO
        // Output registers:
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        STATREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
        );
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_b),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        BUFREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre),
            .lz      (dummy_bufreg_lz[0]),
            .z       (buff)
        );
      end
      else
      begin: CGFIFO
        // Output registers:
        if ( pwropt > 1)
        begin: CGSTATFIFO2
          for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
          begin: pwroptGEN1
            mgc_out_reg
            #(
              .rscid   (rscid),
              .width   (1),
              .ph_clk  (ph_clk),
              .ph_en   (ph_en),
              .ph_arst (ph_arst),
              .ph_srst (ph_srst)
            )
            STATREG
            (
              .clk     (clk),
              .en      (en_l_s[eni/8]),
              .arst    (arst),
              .srst    (srst),
              .ld      (1'b1),
              .d       (stat_pre[eni]),
              .lz      (dummy_statreg_lz[eni]),
              .z       (stat[eni])
            );
          end
        end
        else
        begin: CGSTATFIFO
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          STATREG
          (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
          );
        end
        for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
        begin: pwroptGEN2
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (width),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          BUFREG
          (
            .clk     (clk),
            .en      (en_l[eni]),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre[width*eni+:width]),
            .lz      (dummy_bufreg_lz[eni]),
            .z       (buff[width*eni+:width])
          );
        end
      end
    end
    else
    begin: FEED_THRU
      assign vd = vz;
      assign lz = ld;
      assign z = d;
      assign size = ld && !vz;
    end
    endgenerate

endmodule

//------------------------------------------------------------------
//-- PIPE ENTITIES
//------------------------------------------------------------------
/*
 *
 *             _______________________________________________
 * WRITER    |                                               |          READER
 *           |           MGC_PIPE                            |
 *           |           __________________________          |
 *        --<| vdout  --<| vd ---------------  vz<|-----ldin<|---
 *           |           |      FIFO              |          |
 *        ---|>ldout  ---|>ld ---------------- lz |> ---vdin |>--
 *        ---|>dout -----|>d  ---------------- dz |> ----din |>--
 *           |           |________________________|          |
 *           |_______________________________________________|
 */
// two clock pipe
module mgc_pipe (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, size, req_size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer log2_sz = 3; // log2(fifo_sz)
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer pwropt  = 0; // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output [sz_width-1:0]      size;
    input              req_size;


    mgc_out_fifo_wait_core
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz),
        .pwropt   (pwropt)
    )
    FIFO
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (vdin),
        .vz      (ldin),
        .z       (din),
        .size    (size)
    );

endmodule


//------> C:/PROGRA~1/CALYPT~1/CATAPU~1.126/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
         divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
            rmod = {(width_b){1'b0}} - rmod;
         if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2011a.126 Production Release
//  HLS Date:       Wed Aug  8 00:52:07 PDT 2012
// 
//  Generated by:   oh1015@EEWS104A-005
//  Generated date: Thu Apr 28 15:43:24 2016
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    HSVRGB_core
// ------------------------------------------------------------------


module HSVRGB_core (
  clk, arst_n, r_rsc_mgc_in_wire_d, g_rsc_mgc_in_wire_d, b_rsc_mgc_in_wire_d, H_OUT_rsc_mgc_out_stdreg_d,
      S_OUT_rsc_mgc_out_stdreg_d, V_OUT_rsc_mgc_out_stdreg_d, div_mgc_div_a, div_mgc_div_b,
      div_mgc_div_z, div_mgc_div_1_a, div_mgc_div_1_b, div_mgc_div_1_z, div_mgc_div_2_a,
      div_mgc_div_2_b, div_mgc_div_2_z, div_mgc_div_3_a, div_mgc_div_3_b, div_mgc_div_3_z,
      div_mgc_div_4_a, div_mgc_div_4_b, div_mgc_div_4_z, div_mgc_div_5_a, div_mgc_div_5_b,
      div_mgc_div_5_z, div_mgc_div_6_a, div_mgc_div_6_b, div_mgc_div_6_z, div_mgc_div_7_a,
      div_mgc_div_7_b, div_mgc_div_7_z, div_mgc_div_8_a, div_mgc_div_8_b, div_mgc_div_8_z,
      div_mgc_div_9_a, div_mgc_div_9_b, div_mgc_div_9_z, div_mgc_div_10_a, div_mgc_div_10_b,
      div_mgc_div_10_z, div_mgc_div_11_a, div_mgc_div_11_b, div_mgc_div_11_z, div_mgc_div_12_a,
      div_mgc_div_12_b, div_mgc_div_12_z, div_mgc_div_13_a, div_mgc_div_13_b, div_mgc_div_13_z,
      div_mgc_div_14_a, div_mgc_div_14_b, div_mgc_div_14_z, div_mgc_div_15_a, div_mgc_div_15_b,
      div_mgc_div_15_z_oreg, div_mgc_div_16_a, div_mgc_div_16_b, div_mgc_div_16_z_oreg
);
  input clk;
  input arst_n;
  input [9:0] r_rsc_mgc_in_wire_d;
  input [9:0] g_rsc_mgc_in_wire_d;
  input [9:0] b_rsc_mgc_in_wire_d;
  output [9:0] H_OUT_rsc_mgc_out_stdreg_d;
  reg [9:0] H_OUT_rsc_mgc_out_stdreg_d;
  output [9:0] S_OUT_rsc_mgc_out_stdreg_d;
  reg [9:0] S_OUT_rsc_mgc_out_stdreg_d;
  output [9:0] V_OUT_rsc_mgc_out_stdreg_d;
  reg [9:0] V_OUT_rsc_mgc_out_stdreg_d;
  output [29:0] div_mgc_div_a;
  output [20:0] div_mgc_div_b;
  input [29:0] div_mgc_div_z;
  output [29:0] div_mgc_div_1_a;
  output [20:0] div_mgc_div_1_b;
  input [29:0] div_mgc_div_1_z;
  output [29:0] div_mgc_div_2_a;
  output [20:0] div_mgc_div_2_b;
  input [29:0] div_mgc_div_2_z;
  output [29:0] div_mgc_div_3_a;
  output [20:0] div_mgc_div_3_b;
  input [29:0] div_mgc_div_3_z;
  output [29:0] div_mgc_div_4_a;
  output [20:0] div_mgc_div_4_b;
  input [29:0] div_mgc_div_4_z;
  output [29:0] div_mgc_div_5_a;
  output [20:0] div_mgc_div_5_b;
  input [29:0] div_mgc_div_5_z;
  output [29:0] div_mgc_div_6_a;
  output [20:0] div_mgc_div_6_b;
  input [29:0] div_mgc_div_6_z;
  output [29:0] div_mgc_div_7_a;
  output [20:0] div_mgc_div_7_b;
  input [29:0] div_mgc_div_7_z;
  output [29:0] div_mgc_div_8_a;
  output [20:0] div_mgc_div_8_b;
  input [29:0] div_mgc_div_8_z;
  output [29:0] div_mgc_div_9_a;
  output [20:0] div_mgc_div_9_b;
  input [29:0] div_mgc_div_9_z;
  output [29:0] div_mgc_div_10_a;
  output [20:0] div_mgc_div_10_b;
  input [29:0] div_mgc_div_10_z;
  output [29:0] div_mgc_div_11_a;
  output [20:0] div_mgc_div_11_b;
  input [29:0] div_mgc_div_11_z;
  output [29:0] div_mgc_div_12_a;
  output [20:0] div_mgc_div_12_b;
  input [29:0] div_mgc_div_12_z;
  output [29:0] div_mgc_div_13_a;
  output [20:0] div_mgc_div_13_b;
  input [29:0] div_mgc_div_13_z;
  output [29:0] div_mgc_div_14_a;
  output [20:0] div_mgc_div_14_b;
  input [29:0] div_mgc_div_14_z;
  output [19:0] div_mgc_div_15_a;
  output [9:0] div_mgc_div_15_b;
  input [19:0] div_mgc_div_15_z_oreg;
  output [19:0] div_mgc_div_16_a;
  output [9:0] div_mgc_div_16_b;
  input [19:0] div_mgc_div_16_z_oreg;


  // Interconnect Declarations
  wire [2:0] else_7_if_1_acc_tmp;
  wire [3:0] nl_else_7_if_1_acc_tmp;
  wire [2:0] else_7_else_1_if_acc_tmp;
  wire [3:0] nl_else_7_else_1_if_acc_tmp;
  wire [2:0] else_7_else_1_else_acc_tmp;
  wire [3:0] nl_else_7_else_1_else_acc_tmp;
  wire else_7_else_1_equal_tmp;
  wire else_7_equal_tmp;
  wire [9:0] mux1h_38_tmp;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_74;
  wire and_dcpl_76;
  wire and_dcpl_98;
  wire and_dcpl_136;
  wire and_dcpl_160;
  wire or_tmp_1;
  wire and_dcpl_200;
  wire and_dcpl_201;
  wire and_dcpl_241;
  wire and_dcpl_243;
  wire and_dcpl_261;
  wire and_dcpl_293;
  wire and_dcpl_313;
  wire and_dcpl_348;
  wire and_dcpl_388;
  wire and_dcpl_408;
  wire and_dcpl_440;
  wire and_dcpl_460;
  wire or_tmp_3;
  wire or_tmp_11;
  wire or_tmp_79;
  wire and_dcpl_503;
  wire and_dcpl_504;
  wire and_dcpl_506;
  wire and_dcpl_510;
  wire and_dcpl_515;
  wire and_dcpl_518;
  wire and_dcpl_520;
  wire and_dcpl_521;
  wire and_dcpl_531;
  wire and_dcpl_554;
  wire and_dcpl_555;
  wire and_dcpl_556;
  wire and_dcpl_560;
  wire and_dcpl_562;
  wire and_dcpl_574;
  wire and_dcpl_575;
  wire and_dcpl_588;
  wire and_dcpl_589;
  wire or_dcpl_462;
  wire and_dcpl_626;
  wire and_dcpl_627;
  wire and_dcpl_628;
  wire and_dcpl_630;
  wire and_dcpl_636;
  wire and_dcpl_646;
  wire and_dcpl_647;
  wire and_dcpl_661;
  wire and_dcpl_698;
  wire and_dcpl_699;
  wire and_dcpl_702;
  wire and_dcpl_704;
  wire or_tmp_115;
  wire or_tmp_116;
  wire or_tmp_118;
  wire and_dcpl_709;
  wire or_tmp_123;
  wire mux_tmp_35;
  wire and_dcpl_714;
  wire or_tmp_126;
  wire or_tmp_128;
  wire or_tmp_130;
  wire and_tmp_1;
  wire and_tmp_4;
  wire or_tmp_160;
  wire mux_tmp_46;
  wire and_tmp_9;
  wire nor_tmp_10;
  wire and_tmp_12;
  wire or_tmp_199;
  wire mux_tmp_57;
  wire or_tmp_205;
  wire and_tmp_17;
  wire and_tmp_20;
  wire or_tmp_238;
  wire mux_tmp_68;
  wire and_tmp_25;
  wire nor_tmp_16;
  wire and_tmp_28;
  wire or_tmp_273;
  wire mux_tmp_81;
  wire or_tmp_279;
  wire or_tmp_284;
  wire mux_tmp_84;
  wire or_tmp_295;
  wire mux_tmp_87;
  wire and_dcpl_888;
  wire and_dcpl_889;
  wire and_dcpl_890;
  wire and_dcpl_896;
  wire or_tmp_322;
  wire and_tmp_35;
  wire mux_tmp_99;
  wire or_tmp_330;
  wire and_tmp_37;
  wire and_tmp_40;
  wire or_tmp_363;
  wire mux_tmp_106;
  wire or_tmp_369;
  wire and_tmp_46;
  wire and_tmp_49;
  wire or_tmp_402;
  wire mux_tmp_113;
  wire or_tmp_408;
  wire and_tmp_55;
  wire and_tmp_58;
  wire or_tmp_441;
  wire mux_tmp_120;
  wire or_tmp_447;
  wire and_tmp_64;
  wire and_tmp_67;
  wire nor_tmp_22;
  wire mux_tmp_127;
  wire or_tmp_484;
  wire or_tmp_489;
  wire mux_tmp_129;
  wire or_tmp_500;
  wire mux_tmp_131;
  wire and_dcpl_1118;
  wire and_dcpl_1119;
  wire and_dcpl_1120;
  wire and_dcpl_1126;
  wire or_tmp_527;
  wire and_tmp_75;
  wire mux_tmp_140;
  wire and_tmp_77;
  wire and_tmp_80;
  wire or_tmp_568;
  wire mux_tmp_147;
  wire or_tmp_574;
  wire and_tmp_86;
  wire and_tmp_89;
  wire or_tmp_607;
  wire mux_tmp_154;
  wire or_tmp_613;
  wire and_tmp_95;
  wire and_tmp_98;
  wire or_tmp_646;
  wire mux_tmp_161;
  wire or_tmp_652;
  wire and_tmp_104;
  wire and_tmp_107;
  wire nor_tmp_24;
  wire mux_tmp_168;
  wire or_tmp_689;
  wire or_tmp_694;
  wire mux_tmp_170;
  wire or_tmp_705;
  wire mux_tmp_172;
  wire not_tmp_349;
  wire or_dcpl_790;
  wire or_dcpl_792;
  wire and_dcpl_1348;
  wire and_dcpl_1350;
  wire and_dcpl_1352;
  wire and_dcpl_1354;
  wire or_dcpl_801;
  wire or_dcpl_803;
  wire or_dcpl_805;
  wire or_dcpl_807;
  wire and_tmp_116;
  reg unequal_tmp_1;
  reg else_7_equal_svs;
  reg [10:0] else_7_acc_1_psp_sg1_sva;
  reg else_7_if_div_2cyc;
  reg [17:0] s_sg1_1_sva_2_duc;
  reg [2:0] else_7_if_1_div_5cyc;
  reg [17:0] h_4_sva_duc;
  reg [2:0] else_7_else_1_if_div_5cyc;
  reg [17:0] h_6_sva_duc;
  reg [2:0] else_7_else_1_else_div_5cyc;
  reg [17:0] h_5_sva_duc;
  reg else_7_else_1_equal_svs_1;
  reg else_7_else_1_equal_svs_2;
  reg else_7_else_1_equal_svs_3;
  reg else_7_else_1_equal_svs_4;
  reg else_7_else_1_equal_svs_5;
  reg unequal_tmp_2;
  reg unequal_tmp_3;
  reg unequal_tmp_4;
  reg unequal_tmp_5;
  reg unequal_tmp_6;
  reg unequal_tmp_8;
  reg unequal_tmp_9;
  reg else_7_equal_svs_2;
  reg else_7_equal_svs_3;
  reg else_7_equal_svs_4;
  reg else_7_equal_svs_5;
  reg else_7_and_5_itm_1;
  reg else_7_and_5_itm_2;
  reg else_7_and_5_itm_3;
  reg else_7_and_5_itm_4;
  reg else_7_and_5_itm_5;
  reg [9:0] acc_4_itm_1;
  wire [10:0] nl_acc_4_itm_1;
  reg [9:0] acc_4_itm_2;
  reg [8:0] acc_5_itm_1;
  wire [9:0] nl_acc_5_itm_1;
  reg [8:0] acc_5_itm_2;
  reg [8:0] acc_5_itm_3;
  reg [8:0] acc_5_itm_4;
  reg [8:0] acc_5_itm_5;
  reg [9:0] acc_2_psp_sva_st_1;
  reg else_7_if_div_2cyc_st_1;
  reg [9:0] acc_2_psp_sva_st_2;
  reg [9:0] acc_2_psp_sva_st_3;
  reg [9:0] max_sg1_lpi_dfm_3_st_2;
  reg [9:0] max_sg1_lpi_dfm_3_st_3;
  reg else_7_if_div_2cyc_st_2;
  reg else_7_if_div_2cyc_st_3;
  reg [9:0] acc_2_psp_sva_st_4;
  reg else_7_equal_svs_st_1;
  reg else_7_equal_svs_st_2;
  reg else_7_equal_svs_st_3;
  reg else_7_equal_svs_st_4;
  reg [2:0] else_7_if_1_div_5cyc_st_1;
  reg [2:0] else_7_if_1_div_5cyc_st_2;
  reg [2:0] else_7_if_1_div_5cyc_st_3;
  reg [2:0] else_7_if_1_div_5cyc_st_4;
  reg [9:0] acc_2_psp_sva_st_5;
  reg else_7_equal_svs_st_5;
  reg [2:0] else_7_if_1_div_5cyc_st_5;
  reg else_7_else_1_equal_svs_st_1;
  reg else_7_else_1_equal_svs_st_2;
  reg else_7_else_1_equal_svs_st_3;
  reg else_7_else_1_equal_svs_st_4;
  reg [2:0] else_7_else_1_if_div_5cyc_st_1;
  reg [2:0] else_7_else_1_if_div_5cyc_st_2;
  reg [2:0] else_7_else_1_if_div_5cyc_st_3;
  reg [2:0] else_7_else_1_if_div_5cyc_st_4;
  reg else_7_else_1_equal_svs_st_5;
  reg [2:0] else_7_else_1_if_div_5cyc_st_5;
  reg [2:0] else_7_else_1_else_div_5cyc_st_1;
  reg [2:0] else_7_else_1_else_div_5cyc_st_2;
  reg [2:0] else_7_else_1_else_div_5cyc_st_3;
  reg [2:0] else_7_else_1_else_div_5cyc_st_4;
  reg [2:0] else_7_else_1_else_div_5cyc_st_5;
  reg main_stage_0_2;
  reg main_stage_0_3;
  reg main_stage_0_4;
  reg main_stage_0_5;
  reg main_stage_0_6;
  reg [9:0] else_7_if_conc_1_tmp_mut_sg1;
  reg [9:0] else_7_if_conc_1_tmp_mut_1_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_5_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_6_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_7_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_8_sg1;
  reg [9:0] mut_15_sg1;
  reg [9:0] mut_16_sg1;
  reg [9:0] mut_17_sg1;
  reg [9:0] mut_18_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_5_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_6_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_7_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_8_sg1;
  reg [9:0] mut_19_sg1;
  reg [9:0] mut_20_sg1;
  reg [9:0] mut_21_sg1;
  reg [9:0] mut_22_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_9_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_10_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_11_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_12_sg1;
  reg [9:0] mut_23_sg1;
  reg [9:0] mut_24_sg1;
  reg [9:0] mut_25_sg1;
  reg [9:0] mut_26_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_13_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_14_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_15_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_16_sg1;
  reg [9:0] mut_27_sg1;
  reg [9:0] mut_28_sg1;
  reg [9:0] mut_29_sg1;
  reg [9:0] mut_30_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_17_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_18_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_19_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_20_sg1;
  reg [9:0] mut_31_sg1;
  reg [9:0] mut_32_sg1;
  reg [9:0] mut_33_sg1;
  reg [9:0] mut_34_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_21_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_22_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_23_sg1;
  reg [9:0] else_7_else_1_else_conc_1_tmp_mut_24_sg1;
  reg [9:0] mut_35_sg1;
  reg [9:0] mut_36_sg1;
  reg [9:0] mut_37_sg1;
  reg [9:0] mut_38_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_5_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_6_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_7_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_8_sg1;
  reg [9:0] mut_39_sg1;
  reg [9:0] mut_40_sg1;
  reg [9:0] mut_41_sg1;
  reg [9:0] mut_42_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_9_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_10_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_11_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_12_sg1;
  reg [9:0] mut_43_sg1;
  reg [9:0] mut_44_sg1;
  reg [9:0] mut_45_sg1;
  reg [9:0] mut_46_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_13_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_14_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_15_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_16_sg1;
  reg [9:0] mut_47_sg1;
  reg [9:0] mut_48_sg1;
  reg [9:0] mut_49_sg1;
  reg [9:0] mut_50_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_17_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_18_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_19_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_20_sg1;
  reg [9:0] mut_51_sg1;
  reg [9:0] mut_52_sg1;
  reg [9:0] mut_53_sg1;
  reg [9:0] mut_54_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_21_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_22_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_23_sg1;
  reg [9:0] else_7_else_1_if_conc_1_tmp_mut_24_sg1;
  reg [9:0] mut_55_sg1;
  reg [9:0] mut_56_sg1;
  reg [9:0] mut_57_sg1;
  reg [9:0] mut_58_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_9_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_10_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_11_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_12_sg1;
  reg [9:0] mut_59_sg1;
  reg [9:0] mut_60_sg1;
  reg [9:0] mut_61_sg1;
  reg [9:0] mut_62_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_13_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_14_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_15_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_16_sg1;
  reg [9:0] mut_63_sg1;
  reg [9:0] mut_64_sg1;
  reg [9:0] mut_65_sg1;
  reg [9:0] mut_66_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_17_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_18_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_19_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_20_sg1;
  reg [9:0] mut_67_sg1;
  reg [9:0] mut_68_sg1;
  reg [9:0] mut_69_sg1;
  reg [9:0] mut_70_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_21_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_22_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_23_sg1;
  reg [9:0] else_7_if_1_conc_1_tmp_mut_24_sg1;
  reg [9:0] mut_71_sg1;
  reg [9:0] mut_72_sg1;
  reg [9:0] mut_73_sg1;
  reg [9:0] mut_74_sg1;
  wire and_588_cse;
  wire and_590_cse;
  wire and_592_cse;
  wire and_594_cse;
  wire and_596_cse;
  wire and_660_cse;
  wire and_662_cse;
  wire and_664_cse;
  wire and_666_cse;
  wire and_668_cse;
  wire [5:0] h_4_lpi_dfm_1_sg2_1;
  wire h_4_lpi_dfm_1_sg1_1;
  wire [10:0] h_4_lpi_dfm_4;
  wire or_489_cse;
  wire and_1892_cse;
  wire and_713_cse;
  wire and_718_cse;
  wire and_723_cse;
  wire or_646_cse;
  wire and_764_cse;
  wire and_769_cse;
  wire and_810_cse;
  wire and_815_cse;
  wire and_856_cse;
  wire and_861_cse;
  wire and_902_cse;
  wire and_907_cse;
  wire and_945_cse;
  wire and_952_cse;
  wire and_1000_cse;
  wire and_1007_cse;
  wire and_1055_cse;
  wire and_1062_cse;
  wire and_1110_cse;
  wire and_1117_cse;
  wire and_1165_cse;
  wire and_1172_cse;
  wire and_1215_cse;
  wire and_1222_cse;
  wire and_1270_cse;
  wire and_1277_cse;
  wire and_1325_cse;
  wire and_1332_cse;
  wire and_1380_cse;
  wire and_1387_cse;
  wire and_1435_cse;
  wire and_1442_cse;
  wire and_1483_cse;
  reg [9:0] reg_div_mgc_div_16_b_cse;
  reg [9:0] reg_div_mgc_div_15_b_cse;
  wire nand_11_cse;
  wire or_661_cse;
  wire or_663_cse;
  wire or_718_cse;
  wire or_720_cse;
  wire or_775_cse;
  wire or_777_cse;
  wire nand_22_cse;
  wire nand_23_cse;
  wire or_885_cse;
  wire and_504_cse;
  wire or_946_cse;
  wire or_954_cse;
  wire or_956_cse;
  wire or_1011_cse;
  wire or_1013_cse;
  wire or_1068_cse;
  wire or_1070_cse;
  wire nand_34_cse;
  wire nand_35_cse;
  wire or_1180_cse;
  wire or_1241_cse;
  wire or_1249_cse;
  wire or_1251_cse;
  wire or_1306_cse;
  wire or_1308_cse;
  wire or_1363_cse;
  wire or_1365_cse;
  wire or_1420_cse;
  wire or_1422_cse;
  wire or_1475_cse;
  reg [9:0] reg_div_mgc_div_11_b_tmp;
  reg [9:0] reg_div_mgc_div_11_a_tmp;
  reg [9:0] reg_div_mgc_div_12_b_tmp;
  reg [9:0] reg_div_mgc_div_12_a_tmp;
  reg [9:0] reg_div_mgc_div_13_b_tmp;
  reg [9:0] reg_div_mgc_div_13_a_tmp;
  reg [9:0] reg_div_mgc_div_14_b_tmp;
  reg [9:0] reg_div_mgc_div_14_a_tmp;
  reg [9:0] reg_div_mgc_div_b_tmp;
  reg [9:0] reg_div_mgc_div_a_tmp;
  reg [9:0] reg_div_mgc_div_6_b_tmp;
  reg [9:0] reg_div_mgc_div_6_a_tmp;
  reg [9:0] reg_div_mgc_div_7_b_tmp;
  reg [9:0] reg_div_mgc_div_7_a_tmp;
  reg [9:0] reg_div_mgc_div_8_b_tmp;
  reg [9:0] reg_div_mgc_div_8_a_tmp;
  reg [9:0] reg_div_mgc_div_9_b_tmp;
  reg [9:0] reg_div_mgc_div_9_a_tmp;
  reg [9:0] reg_div_mgc_div_10_b_tmp;
  reg [9:0] reg_div_mgc_div_10_a_tmp;
  reg [9:0] reg_div_mgc_div_1_b_tmp;
  reg [9:0] reg_div_mgc_div_1_a_tmp;
  reg [9:0] reg_div_mgc_div_2_b_tmp;
  reg [9:0] reg_div_mgc_div_2_a_tmp;
  reg [9:0] reg_div_mgc_div_3_b_tmp;
  reg [9:0] reg_div_mgc_div_3_a_tmp;
  reg [9:0] reg_div_mgc_div_4_b_tmp;
  reg [9:0] reg_div_mgc_div_4_a_tmp;
  reg [9:0] reg_div_mgc_div_5_b_tmp;
  reg [9:0] reg_div_mgc_div_5_a_tmp;
  wire and_759_cse;
  wire and_805_cse;
  wire and_851_cse;
  wire and_897_cse;
  wire and_938_cse;
  wire and_994_cse;
  wire and_1049_cse;
  wire and_1104_cse;
  wire and_1159_cse;
  wire and_1208_cse;
  wire and_1264_cse;
  wire and_1319_cse;
  wire and_1374_cse;
  wire and_1429_cse;
  reg [9:0] reg_max_sg1_lpi_dfm_3_st_1_cse;
  wire and_304_cse;
  wire and_146_cse;
  wire and_356_cse;
  wire and_208_cse;
  wire mux_143_cse;
  wire mux_187_cse;
  wire mux_228_cse;
  wire and_730_cse;
  wire mux_95_cse;
  wire and_776_cse;
  wire mux_106_cse;
  wire and_822_cse;
  wire mux_117_cse;
  wire and_868_cse;
  wire mux_128_cse;
  wire and_913_cse;
  wire and_960_cse;
  wire mux_157_cse;
  wire and_1015_cse;
  wire mux_164_cse;
  wire and_1070_cse;
  wire mux_171_cse;
  wire and_1125_cse;
  wire mux_178_cse;
  wire and_1179_cse;
  wire and_1230_cse;
  wire mux_198_cse;
  wire and_1285_cse;
  wire mux_205_cse;
  wire and_1340_cse;
  wire mux_212_cse;
  wire and_1395_cse;
  wire mux_219_cse;
  wire and_1449_cse;
  wire mux_145_cse;
  wire mux_188_cse;
  wire mux_229_cse;
  wire [17:0] else_7_acc_1_itm;
  wire [18:0] nl_else_7_acc_1_itm;
  wire [10:0] acc_itm;
  wire [11:0] nl_acc_itm;
  wire [10:0] else_7_acc_1_psp_sg1_sva_1;
  wire [17:0] h_4_sva_duc_mx0;
  wire [6:0] h_4_sva_1_sg1;
  wire [7:0] nl_h_4_sva_1_sg1;
  wire [17:0] h_5_sva_duc_mx0;
  wire else_7_nor_ssc;
  wire [3:0] h_1_sg1_lpi_dfm_1;
  wire [2:0] acc_imod;
  wire [3:0] nl_acc_imod;
  wire [2:0] else_7_if_1_acc_idiv;
  wire [3:0] nl_else_7_if_1_acc_idiv;
  wire [9:0] g_1_lpi_dfm;
  wire [9:0] b_1_lpi_dfm;
  wire [2:0] acc_imod_1;
  wire [3:0] nl_acc_imod_1;
  wire [2:0] else_7_else_1_if_acc_idiv;
  wire [3:0] nl_else_7_else_1_if_acc_idiv;
  wire [9:0] r_1_lpi_dfm;
  wire [2:0] acc_imod_2;
  wire [3:0] nl_acc_imod_2;
  wire [2:0] else_7_else_1_else_acc_idiv;
  wire [3:0] nl_else_7_else_1_else_acc_idiv;
  wire unequal_tmp_10;
  wire or_cse;
  wire [11:0] if_if_acc_itm;
  wire [12:0] nl_if_if_acc_itm;
  wire [11:0] else_1_if_acc_itm;
  wire [12:0] nl_else_1_if_acc_itm;
  wire [11:0] if_3_if_acc_itm;
  wire [12:0] nl_if_3_if_acc_itm;
  wire [11:0] else_5_if_acc_itm;
  wire [12:0] nl_else_5_if_acc_itm;
  wire [10:0] else_7_if_1_acc_1_itm;
  wire [11:0] nl_else_7_if_1_acc_1_itm;
  wire [10:0] else_7_else_1_if_acc_2_itm;
  wire [11:0] nl_else_7_else_1_if_acc_2_itm;
  wire [10:0] else_7_else_1_else_acc_2_itm;
  wire [11:0] nl_else_7_else_1_else_acc_2_itm;
  wire [11:0] if_3_acc_1_itm;
  wire [12:0] nl_if_3_acc_1_itm;
  wire [11:0] if_acc_1_itm;
  wire [12:0] nl_if_acc_1_itm;
  wire [17:0] mul_1_itm;
  wire [35:0] nl_mul_1_itm;
  wire [13:0] mul_itm;
  wire [27:0] nl_mul_itm;

  wire[0:0] mux_88_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] mux_224_nl;
  wire[6:0] mux1h_3_nl;
  wire[5:0] mux1h_6_nl;
  wire[9:0] mux1h_39_nl;
  wire[17:0] mux1h_40_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_226_nl;

  // Interconnect Declarations for Component Instantiations 
  assign and_1892_cse = (~((acc_2_psp_sva_st_5[7]) | (acc_2_psp_sva_st_5[6]) | (acc_2_psp_sva_st_5[5])))
      & (~((acc_2_psp_sva_st_5[4]) | (acc_2_psp_sva_st_5[3]))) & (~((acc_2_psp_sva_st_5[2])
      | (acc_2_psp_sva_st_5[1]) | (acc_2_psp_sva_st_5[0]))) & (~((acc_2_psp_sva_st_5[9])
      | (acc_2_psp_sva_st_5[8])));
  assign or_489_cse = (acc_2_psp_sva_st_5[7]) | (acc_2_psp_sva_st_5[6]) | (acc_2_psp_sva_st_5[5])
      | (acc_2_psp_sva_st_5[4]) | (acc_2_psp_sva_st_5[3]) | (acc_2_psp_sva_st_5[2])
      | (acc_2_psp_sva_st_5[1]) | (acc_2_psp_sva_st_5[0]) | (acc_2_psp_sva_st_5[9])
      | (acc_2_psp_sva_st_5[8]);
  assign or_646_cse = (acc_itm[1]) | (acc_itm[2]) | (acc_itm[3]) | (acc_itm[4]) |
      (acc_itm[5]) | (acc_itm[6]) | (acc_itm[7]) | (acc_itm[8]) | (acc_itm[9]) |
      (acc_itm[10]);
  assign and_713_cse = or_646_cse & and_dcpl_699 & and_dcpl_698;
  assign mux_88_nl = MUX_s_1_2_2({(~ or_tmp_118) , or_tmp_116}, or_tmp_115);
  assign and_718_cse = (mux_88_nl) & and_dcpl_704 & and_dcpl_702;
  assign mux_91_nl = MUX_s_1_2_2({(nand_11_cse & mux_tmp_35) , mux_tmp_35}, or_tmp_115);
  assign and_723_cse = (mux_91_nl) & and_dcpl_709 & and_dcpl_200;
  assign div_mgc_div_11_b = {1'b0, {reg_div_mgc_div_11_b_tmp , 10'b0}};
  assign div_mgc_div_11_a = {reg_div_mgc_div_11_a_tmp , 20'b0};
  assign mux_100_nl = MUX_s_1_2_2({(~ or_tmp_118) , or_tmp_116}, or_tmp_160);
  assign and_764_cse = (mux_100_nl) & and_dcpl_704 & (else_7_if_1_div_5cyc_st_1[0])
      & (~ (else_7_if_1_div_5cyc_st_1[1]));
  assign mux_102_nl = MUX_s_1_2_2({(nand_11_cse & mux_tmp_46) , mux_tmp_46}, or_tmp_160);
  assign and_769_cse = (mux_102_nl) & and_dcpl_709 & (~ (else_7_if_1_div_5cyc_st_2[1]))
      & (else_7_if_1_div_5cyc_st_2[0]);
  assign and_759_cse = or_646_cse & and_dcpl_699 & (~ (else_7_if_1_acc_tmp[1])) &
      (else_7_if_1_acc_tmp[0]);
  assign div_mgc_div_12_b = {1'b0, {reg_div_mgc_div_12_b_tmp , 10'b0}};
  assign div_mgc_div_12_a = {reg_div_mgc_div_12_a_tmp , 20'b0};
  assign mux_111_nl = MUX_s_1_2_2({(~ or_tmp_118) , or_tmp_116}, or_tmp_199);
  assign and_810_cse = (mux_111_nl) & and_dcpl_704 & (~ (else_7_if_1_div_5cyc_st_1[0]))
      & (else_7_if_1_div_5cyc_st_1[1]);
  assign mux_113_nl = MUX_s_1_2_2({(nand_11_cse & mux_tmp_57) , mux_tmp_57}, or_tmp_199);
  assign and_815_cse = (mux_113_nl) & and_dcpl_709 & (else_7_if_1_div_5cyc_st_2[1])
      & (~ (else_7_if_1_div_5cyc_st_2[0]));
  assign and_805_cse = or_646_cse & and_dcpl_699 & (else_7_if_1_acc_tmp[1]) & (~
      (else_7_if_1_acc_tmp[0]));
  assign div_mgc_div_13_b = {1'b0, {reg_div_mgc_div_13_b_tmp , 10'b0}};
  assign div_mgc_div_13_a = {reg_div_mgc_div_13_a_tmp , 20'b0};
  assign mux_122_nl = MUX_s_1_2_2({(~ or_tmp_118) , or_tmp_116}, or_tmp_238);
  assign and_856_cse = (mux_122_nl) & and_dcpl_704 & (else_7_if_1_div_5cyc_st_1[0])
      & (else_7_if_1_div_5cyc_st_1[1]);
  assign mux_124_nl = MUX_s_1_2_2({(nand_11_cse & mux_tmp_68) , mux_tmp_68}, or_tmp_238);
  assign and_861_cse = (mux_124_nl) & and_dcpl_709 & (else_7_if_1_div_5cyc_st_2[1])
      & (else_7_if_1_div_5cyc_st_2[0]);
  assign and_851_cse = or_646_cse & and_dcpl_699 & (else_7_if_1_acc_tmp[1]) & (else_7_if_1_acc_tmp[0]);
  assign div_mgc_div_14_b = {1'b0, {reg_div_mgc_div_14_b_tmp , 10'b0}};
  assign div_mgc_div_14_a = {reg_div_mgc_div_14_a_tmp , 20'b0};
  assign mux_133_nl = MUX_s_1_2_2({or_tmp_116 , (~ or_tmp_118)}, else_7_if_1_acc_tmp[2]);
  assign mux_134_nl = MUX_s_1_2_2({(mux_133_nl) , or_tmp_116}, or_tmp_273);
  assign and_902_cse = (mux_134_nl) & and_dcpl_348 & (else_7_if_1_div_5cyc_st_1[2])
      & and_dcpl_702;
  assign mux_137_nl = MUX_s_1_2_2({mux_tmp_81 , (nand_11_cse & mux_tmp_81)}, else_7_if_1_acc_tmp[2]);
  assign mux_138_nl = MUX_s_1_2_2({(mux_137_nl) , mux_tmp_81}, or_tmp_273);
  assign and_907_cse = (mux_138_nl) & and_dcpl_201 & (else_7_if_1_div_5cyc_st_2[2])
      & and_dcpl_200;
  assign and_897_cse = or_646_cse & else_7_equal_tmp & (else_7_if_1_acc_tmp[2]) &
      and_dcpl_698;
  assign div_mgc_div_b = {1'b0, {reg_div_mgc_div_b_tmp , 10'b0}};
  assign div_mgc_div_a = {reg_div_mgc_div_a_tmp , 20'b0};
  assign mux_153_nl = MUX_s_1_2_2({and_tmp_35 , or_tmp_116}, or_tmp_322);
  assign and_945_cse = (mux_153_nl) & and_dcpl_896 & and_dcpl_388 & (~ (else_7_else_1_if_div_5cyc_st_1[0]));
  assign mux_155_nl = MUX_s_1_2_2({(or_946_cse & mux_tmp_99) , mux_tmp_99}, or_tmp_322);
  assign and_952_cse = (mux_155_nl) & and_304_cse & and_dcpl_241 & (~ (else_7_else_1_if_div_5cyc_st_2[0]));
  assign and_938_cse = or_646_cse & and_dcpl_890 & and_dcpl_888;
  assign div_mgc_div_6_b = {1'b0, {reg_div_mgc_div_6_b_tmp , 10'b0}};
  assign div_mgc_div_6_a = {reg_div_mgc_div_6_a_tmp , 20'b0};
  assign mux_160_nl = MUX_s_1_2_2({and_tmp_35 , or_tmp_116}, or_tmp_363);
  assign and_1000_cse = (mux_160_nl) & and_dcpl_896 & and_dcpl_388 & (else_7_else_1_if_div_5cyc_st_1[0]);
  assign mux_162_nl = MUX_s_1_2_2({(or_946_cse & mux_tmp_106) , mux_tmp_106}, or_tmp_363);
  assign and_1007_cse = (mux_162_nl) & and_304_cse & and_dcpl_241 & (else_7_else_1_if_div_5cyc_st_2[0]);
  assign and_994_cse = or_646_cse & and_dcpl_890 & (~ (else_7_else_1_if_acc_tmp[1]))
      & (else_7_else_1_if_acc_tmp[0]);
  assign div_mgc_div_7_b = {1'b0, {reg_div_mgc_div_7_b_tmp , 10'b0}};
  assign div_mgc_div_7_a = {reg_div_mgc_div_7_a_tmp , 20'b0};
  assign mux_167_nl = MUX_s_1_2_2({and_tmp_35 , or_tmp_116}, or_tmp_402);
  assign and_1055_cse = (mux_167_nl) & and_dcpl_896 & and_dcpl_408 & (~ (else_7_else_1_if_div_5cyc_st_1[0]));
  assign mux_169_nl = MUX_s_1_2_2({(or_946_cse & mux_tmp_113) , mux_tmp_113}, or_tmp_402);
  assign and_1062_cse = (mux_169_nl) & and_304_cse & and_dcpl_261 & (~ (else_7_else_1_if_div_5cyc_st_2[0]));
  assign and_1049_cse = or_646_cse & and_dcpl_890 & (else_7_else_1_if_acc_tmp[1])
      & (~ (else_7_else_1_if_acc_tmp[0]));
  assign div_mgc_div_8_b = {1'b0, {reg_div_mgc_div_8_b_tmp , 10'b0}};
  assign div_mgc_div_8_a = {reg_div_mgc_div_8_a_tmp , 20'b0};
  assign mux_174_nl = MUX_s_1_2_2({and_tmp_35 , or_tmp_116}, or_tmp_441);
  assign and_1110_cse = (mux_174_nl) & and_dcpl_896 & and_dcpl_408 & (else_7_else_1_if_div_5cyc_st_1[0]);
  assign mux_176_nl = MUX_s_1_2_2({(or_946_cse & mux_tmp_120) , mux_tmp_120}, or_tmp_441);
  assign and_1117_cse = (mux_176_nl) & and_304_cse & and_dcpl_261 & (else_7_else_1_if_div_5cyc_st_2[0]);
  assign and_1104_cse = or_646_cse & and_dcpl_890 & (else_7_else_1_if_acc_tmp[1])
      & (else_7_else_1_if_acc_tmp[0]);
  assign div_mgc_div_9_b = {1'b0, {reg_div_mgc_div_9_b_tmp , 10'b0}};
  assign div_mgc_div_9_a = {reg_div_mgc_div_9_a_tmp , 20'b0};
  assign mux_181_nl = MUX_s_1_2_2({or_tmp_116 , and_tmp_35}, nor_tmp_22);
  assign and_1165_cse = (mux_181_nl) & and_dcpl_896 & (else_7_else_1_if_div_5cyc_st_1[2])
      & (~ (else_7_else_1_if_div_5cyc_st_1[1])) & (~ (else_7_else_1_if_div_5cyc_st_1[0]));
  assign mux_183_nl = MUX_s_1_2_2({mux_tmp_127 , (or_946_cse & mux_tmp_127)}, nor_tmp_22);
  assign and_1172_cse = (mux_183_nl) & and_304_cse & (else_7_else_1_if_div_5cyc_st_2[2])
      & (~ (else_7_else_1_if_div_5cyc_st_2[1])) & (~ (else_7_else_1_if_div_5cyc_st_2[0]));
  assign and_1159_cse = or_646_cse & and_dcpl_889 & (else_7_else_1_if_acc_tmp[2])
      & and_dcpl_888;
  assign div_mgc_div_10_b = {1'b0, {reg_div_mgc_div_10_b_tmp , 10'b0}};
  assign div_mgc_div_10_a = {reg_div_mgc_div_10_a_tmp , 20'b0};
  assign mux_194_nl = MUX_s_1_2_2({and_tmp_75 , or_tmp_116}, or_tmp_527);
  assign and_1215_cse = (mux_194_nl) & and_dcpl_1126 & and_dcpl_440 & (~ (else_7_else_1_else_div_5cyc_st_1[0]));
  assign mux_196_nl = MUX_s_1_2_2({(or_1241_cse & mux_tmp_140) , mux_tmp_140}, or_tmp_527);
  assign and_1222_cse = (mux_196_nl) & and_356_cse & and_dcpl_293 & (~ (else_7_else_1_else_div_5cyc_st_2[0]));
  assign and_1208_cse = or_646_cse & and_dcpl_1120 & and_dcpl_1118;
  assign div_mgc_div_1_b = {1'b0, {reg_div_mgc_div_1_b_tmp , 10'b0}};
  assign div_mgc_div_1_a = {reg_div_mgc_div_1_a_tmp , 20'b0};
  assign mux_201_nl = MUX_s_1_2_2({and_tmp_75 , or_tmp_116}, or_tmp_568);
  assign and_1270_cse = (mux_201_nl) & and_dcpl_1126 & and_dcpl_440 & (else_7_else_1_else_div_5cyc_st_1[0]);
  assign mux_203_nl = MUX_s_1_2_2({(or_1241_cse & mux_tmp_147) , mux_tmp_147}, or_tmp_568);
  assign and_1277_cse = (mux_203_nl) & and_356_cse & and_dcpl_293 & (else_7_else_1_else_div_5cyc_st_2[0]);
  assign and_1264_cse = or_646_cse & and_dcpl_1120 & (~ (else_7_else_1_else_acc_tmp[1]))
      & (else_7_else_1_else_acc_tmp[0]);
  assign div_mgc_div_2_b = {1'b0, {reg_div_mgc_div_2_b_tmp , 10'b0}};
  assign div_mgc_div_2_a = {reg_div_mgc_div_2_a_tmp , 20'b0};
  assign mux_208_nl = MUX_s_1_2_2({and_tmp_75 , or_tmp_116}, or_tmp_607);
  assign and_1325_cse = (mux_208_nl) & and_dcpl_1126 & and_dcpl_460 & (~ (else_7_else_1_else_div_5cyc_st_1[0]));
  assign mux_210_nl = MUX_s_1_2_2({(or_1241_cse & mux_tmp_154) , mux_tmp_154}, or_tmp_607);
  assign and_1332_cse = (mux_210_nl) & and_356_cse & and_dcpl_313 & (~ (else_7_else_1_else_div_5cyc_st_2[0]));
  assign and_1319_cse = or_646_cse & and_dcpl_1120 & (else_7_else_1_else_acc_tmp[1])
      & (~ (else_7_else_1_else_acc_tmp[0]));
  assign div_mgc_div_3_b = {1'b0, {reg_div_mgc_div_3_b_tmp , 10'b0}};
  assign div_mgc_div_3_a = {reg_div_mgc_div_3_a_tmp , 20'b0};
  assign mux_215_nl = MUX_s_1_2_2({and_tmp_75 , or_tmp_116}, or_tmp_646);
  assign and_1380_cse = (mux_215_nl) & and_dcpl_1126 & and_dcpl_460 & (else_7_else_1_else_div_5cyc_st_1[0]);
  assign mux_217_nl = MUX_s_1_2_2({(or_1241_cse & mux_tmp_161) , mux_tmp_161}, or_tmp_646);
  assign and_1387_cse = (mux_217_nl) & and_356_cse & and_dcpl_313 & (else_7_else_1_else_div_5cyc_st_2[0]);
  assign and_1374_cse = or_646_cse & and_dcpl_1120 & (else_7_else_1_else_acc_tmp[1])
      & (else_7_else_1_else_acc_tmp[0]);
  assign div_mgc_div_4_b = {1'b0, {reg_div_mgc_div_4_b_tmp , 10'b0}};
  assign div_mgc_div_4_a = {reg_div_mgc_div_4_a_tmp , 20'b0};
  assign mux_222_nl = MUX_s_1_2_2({or_tmp_116 , and_tmp_75}, nor_tmp_24);
  assign and_1435_cse = (mux_222_nl) & and_dcpl_1126 & (else_7_else_1_else_div_5cyc_st_1[2])
      & (~ (else_7_else_1_else_div_5cyc_st_1[1])) & (~ (else_7_else_1_else_div_5cyc_st_1[0]));
  assign mux_224_nl = MUX_s_1_2_2({mux_tmp_168 , (or_1241_cse & mux_tmp_168)}, nor_tmp_24);
  assign and_1442_cse = (mux_224_nl) & and_356_cse & (~ (else_7_else_1_else_div_5cyc_st_2[1]))
      & (else_7_else_1_else_div_5cyc_st_2[2]) & (~ (else_7_else_1_else_div_5cyc_st_2[0]));
  assign and_1429_cse = or_646_cse & and_dcpl_1119 & (else_7_else_1_else_acc_tmp[2])
      & and_dcpl_1118;
  assign div_mgc_div_5_b = {1'b0, {reg_div_mgc_div_5_b_tmp , 10'b0}};
  assign div_mgc_div_5_a = {reg_div_mgc_div_5_a_tmp , 20'b0};
  assign and_146_cse = and_dcpl_76 & else_7_else_1_equal_svs_st_3;
  assign and_208_cse = and_dcpl_76 & (~ else_7_else_1_equal_svs_st_3);
  assign and_304_cse = and_dcpl_243 & else_7_else_1_equal_svs_st_2;
  assign and_356_cse = and_dcpl_243 & (~ else_7_else_1_equal_svs_st_2);
  assign and_504_cse = main_stage_0_2 & (~ else_7_equal_svs_st_1);
  assign div_mgc_div_16_b = reg_div_mgc_div_16_b_cse;
  assign div_mgc_div_16_a = {else_7_if_conc_1_tmp_mut_1_sg1 , 10'b0};
  assign div_mgc_div_15_b = reg_div_mgc_div_15_b_cse;
  assign div_mgc_div_15_a = {else_7_if_conc_1_tmp_mut_sg1 , 10'b0};
  assign and_1483_cse = and_dcpl_1354 & and_dcpl_1352 & and_dcpl_1350 & and_dcpl_1348;
  assign or_cse = (acc_itm[10]) | (acc_itm[9]) | (acc_itm[8]) | (acc_itm[7]) | (acc_itm[6])
      | (acc_itm[5]) | (acc_itm[4]) | (acc_itm[3]) | (acc_itm[2]) | (acc_itm[1]);
  assign else_7_acc_1_psp_sg1_sva_1 = MUX_v_11_2_2({(else_7_acc_1_itm[17:7]) , else_7_acc_1_psp_sg1_sva},
      and_1892_cse);
  assign nl_else_7_acc_1_itm = ({(~ h_4_lpi_dfm_1_sg2_1) , (~ h_4_lpi_dfm_1_sg1_1)
      , (~ h_4_lpi_dfm_4)}) + ({(h_4_lpi_dfm_1_sg2_1[1:0]) , h_4_lpi_dfm_1_sg1_1
      , h_4_lpi_dfm_4 , 4'b1});
  assign else_7_acc_1_itm = nl_else_7_acc_1_itm[17:0];
  assign h_4_sva_duc_mx0 = MUX1HOT_v_18_6_2({(div_mgc_div_11_z[17:0]) , (div_mgc_div_12_z[17:0])
      , (div_mgc_div_13_z[17:0]) , (div_mgc_div_14_z[17:0]) , (div_mgc_div_z[17:0])
      , h_4_sva_duc}, {(and_dcpl_504 & and_dcpl_503) , (and_dcpl_504 & and_dcpl_506)
      , (and_dcpl_510 & and_dcpl_503) , (and_dcpl_510 & and_dcpl_506) , (and_dcpl_504
      & and_dcpl_515) , (and_dcpl_518 | (~ else_7_equal_svs_st_5))});
  assign mux1h_3_nl = MUX1HOT_v_7_6_2({(div_mgc_div_6_z[17:11]) , (div_mgc_div_7_z[17:11])
      , (div_mgc_div_8_z[17:11]) , (div_mgc_div_9_z[17:11]) , (div_mgc_div_10_z[17:11])
      , (h_6_sva_duc[17:11])}, {and_588_cse , and_590_cse , and_592_cse , and_594_cse
      , and_596_cse , and_dcpl_574});
  assign nl_h_4_sva_1_sg1 = (mux1h_3_nl) + 7'b1;
  assign h_4_sva_1_sg1 = nl_h_4_sva_1_sg1[6:0];
  assign h_5_sva_duc_mx0 = MUX1HOT_v_18_6_2({(div_mgc_div_1_z[17:0]) , (div_mgc_div_2_z[17:0])
      , (div_mgc_div_3_z[17:0]) , (div_mgc_div_4_z[17:0]) , (div_mgc_div_5_z[17:0])
      , h_5_sva_duc}, {(and_dcpl_628 & and_dcpl_626) , (and_dcpl_628 & and_dcpl_630)
      , (and_dcpl_636 & and_dcpl_626) , (and_dcpl_636 & and_dcpl_630) , (and_dcpl_628
      & (~ (else_7_else_1_else_div_5cyc_st_5[0])) & (else_7_else_1_else_div_5cyc_st_5[2]))
      , (and_dcpl_646 | else_7_equal_svs_st_5 | else_7_else_1_equal_svs_st_5)});
  assign mux1h_6_nl = MUX1HOT_v_6_6_2({(div_mgc_div_1_z[17:12]) , (div_mgc_div_2_z[17:12])
      , (div_mgc_div_3_z[17:12]) , (div_mgc_div_4_z[17:12]) , (div_mgc_div_5_z[17:12])
      , (h_5_sva_duc[17:12])}, {and_660_cse , and_662_cse , and_664_cse , and_666_cse
      , and_668_cse , and_dcpl_646});
  assign h_4_lpi_dfm_1_sg2_1 = MUX1HOT_v_6_3_2({((mux1h_6_nl) + 6'b1) , (h_4_sva_1_sg1[6:1])
      , (h_4_sva_duc_mx0[17:12])}, {else_7_nor_ssc , else_7_and_5_itm_5 , else_7_equal_svs_5});
  assign h_4_lpi_dfm_1_sg1_1 = MUX1HOT_s_1_3_2({(h_5_sva_duc_mx0[11]) , (h_4_sva_1_sg1[0])
      , (h_4_sva_duc_mx0[11])}, {else_7_nor_ssc , else_7_and_5_itm_5 , else_7_equal_svs_5});
  assign h_4_lpi_dfm_4 = MUX1HOT_v_11_8_2({(h_5_sva_duc_mx0[10:0]) , (div_mgc_div_6_z[10:0])
      , (div_mgc_div_7_z[10:0]) , (div_mgc_div_8_z[10:0]) , (div_mgc_div_9_z[10:0])
      , (div_mgc_div_10_z[10:0]) , (h_6_sva_duc[10:0]) , (h_4_sva_duc_mx0[10:0])},
      {else_7_nor_ssc , (and_dcpl_556 & and_dcpl_554 & else_7_and_5_itm_5) , (and_dcpl_560
      & and_dcpl_554 & else_7_and_5_itm_5) , (and_dcpl_556 & and_dcpl_562 & else_7_and_5_itm_5)
      , (and_dcpl_560 & and_dcpl_562 & else_7_and_5_itm_5) , (and_dcpl_556 & (~ (else_7_else_1_if_div_5cyc_st_5[1]))
      & (else_7_else_1_if_div_5cyc_st_5[2]) & else_7_and_5_itm_5) , ((and_dcpl_574
      | else_7_equal_svs_st_5 | (~ else_7_else_1_equal_svs_st_5)) & else_7_and_5_itm_5)
      , else_7_equal_svs_5});
  assign else_7_nor_ssc = ~(else_7_else_1_equal_svs_5 | else_7_equal_svs_5);
  assign h_1_sg1_lpi_dfm_1 = (else_7_acc_1_psp_sg1_sva_1[3:0]) & ({{3{unequal_tmp_6}},
      unequal_tmp_6});
  assign nl_if_if_acc_itm = ({1'b1 , r_rsc_mgc_in_wire_d , 1'b1}) + conv_u2u_11_12({(~
      b_rsc_mgc_in_wire_d) , 1'b1});
  assign if_if_acc_itm = nl_if_if_acc_itm[11:0];
  assign nl_else_1_if_acc_itm = ({1'b1 , g_rsc_mgc_in_wire_d , 1'b1}) + conv_u2u_11_12({(~
      b_rsc_mgc_in_wire_d) , 1'b1});
  assign else_1_if_acc_itm = nl_else_1_if_acc_itm[11:0];
  assign nl_if_3_if_acc_itm = ({1'b1 , b_rsc_mgc_in_wire_d , 1'b1}) + conv_u2u_11_12({(~
      r_rsc_mgc_in_wire_d) , 1'b1});
  assign if_3_if_acc_itm = nl_if_3_if_acc_itm[11:0];
  assign nl_else_5_if_acc_itm = ({1'b1 , b_rsc_mgc_in_wire_d , 1'b1}) + conv_u2u_11_12({(~
      g_rsc_mgc_in_wire_d) , 1'b1});
  assign else_5_if_acc_itm = nl_else_5_if_acc_itm[11:0];
  assign mux1h_38_tmp = MUX1HOT_v_10_3_2({r_rsc_mgc_in_wire_d , b_rsc_mgc_in_wire_d
      , g_rsc_mgc_in_wire_d}, {(~((if_if_acc_itm[11]) | (if_acc_1_itm[11]))) , (((if_if_acc_itm[11])
      & (~ (if_acc_1_itm[11]))) | ((else_1_if_acc_itm[11]) & (if_acc_1_itm[11])))
      , ((~ (else_1_if_acc_itm[11])) & (if_acc_1_itm[11]))});
  assign mux1h_39_nl = MUX1HOT_v_10_3_2({r_rsc_mgc_in_wire_d , b_rsc_mgc_in_wire_d
      , g_rsc_mgc_in_wire_d}, {(~((if_3_if_acc_itm[11]) | (if_3_acc_1_itm[11])))
      , (((if_3_if_acc_itm[11]) & (~ (if_3_acc_1_itm[11]))) | ((else_5_if_acc_itm[11])
      & (if_3_acc_1_itm[11]))) , ((~ (else_5_if_acc_itm[11])) & (if_3_acc_1_itm[11]))});
  assign nl_acc_itm = ({mux1h_38_tmp , 1'b1}) + ({(~ (mux1h_39_nl)) , 1'b1});
  assign acc_itm = nl_acc_itm[10:0];
  assign nl_else_7_if_1_acc_1_itm = ({g_1_lpi_dfm , 1'b1}) + ({(~ b_1_lpi_dfm) ,
      1'b1});
  assign else_7_if_1_acc_1_itm = nl_else_7_if_1_acc_1_itm[10:0];
  assign nl_else_7_if_1_acc_tmp = conv_u2u_1_3(acc_imod[2]) + conv_u2u_2_3(acc_imod[1:0]);
  assign else_7_if_1_acc_tmp = nl_else_7_if_1_acc_tmp[2:0];
  assign nl_acc_imod = conv_s2s_1_3(else_7_if_1_acc_idiv[2]) + conv_u2s_2_3(else_7_if_1_acc_idiv[1:0]);
  assign acc_imod = nl_acc_imod[2:0];
  assign nl_else_7_if_1_acc_idiv = else_7_if_1_div_5cyc + 3'b1;
  assign else_7_if_1_acc_idiv = nl_else_7_if_1_acc_idiv[2:0];
  assign g_1_lpi_dfm = g_rsc_mgc_in_wire_d & ({{9{unequal_tmp_10}}, unequal_tmp_10});
  assign b_1_lpi_dfm = b_rsc_mgc_in_wire_d & ({{9{unequal_tmp_10}}, unequal_tmp_10});
  assign nl_else_7_else_1_if_acc_2_itm = ({b_1_lpi_dfm , 1'b1}) + ({(~ r_1_lpi_dfm)
      , 1'b1});
  assign else_7_else_1_if_acc_2_itm = nl_else_7_else_1_if_acc_2_itm[10:0];
  assign nl_else_7_else_1_if_acc_tmp = conv_u2u_1_3(acc_imod_1[2]) + conv_u2u_2_3(acc_imod_1[1:0]);
  assign else_7_else_1_if_acc_tmp = nl_else_7_else_1_if_acc_tmp[2:0];
  assign nl_acc_imod_1 = conv_s2s_1_3(else_7_else_1_if_acc_idiv[2]) + conv_u2s_2_3(else_7_else_1_if_acc_idiv[1:0]);
  assign acc_imod_1 = nl_acc_imod_1[2:0];
  assign nl_else_7_else_1_if_acc_idiv = else_7_else_1_if_div_5cyc + 3'b1;
  assign else_7_else_1_if_acc_idiv = nl_else_7_else_1_if_acc_idiv[2:0];
  assign r_1_lpi_dfm = r_rsc_mgc_in_wire_d & ({{9{unequal_tmp_10}}, unequal_tmp_10});
  assign nl_else_7_else_1_else_acc_2_itm = ({r_1_lpi_dfm , 1'b1}) + ({(~ g_1_lpi_dfm)
      , 1'b1});
  assign else_7_else_1_else_acc_2_itm = nl_else_7_else_1_else_acc_2_itm[10:0];
  assign nl_else_7_else_1_else_acc_tmp = conv_u2u_1_3(acc_imod_2[2]) + conv_u2u_2_3(acc_imod_2[1:0]);
  assign else_7_else_1_else_acc_tmp = nl_else_7_else_1_else_acc_tmp[2:0];
  assign nl_acc_imod_2 = conv_s2s_1_3(else_7_else_1_else_acc_idiv[2]) + conv_u2s_2_3(else_7_else_1_else_acc_idiv[1:0]);
  assign acc_imod_2 = nl_acc_imod_2[2:0];
  assign nl_else_7_else_1_else_acc_idiv = else_7_else_1_else_div_5cyc + 3'b1;
  assign else_7_else_1_else_acc_idiv = nl_else_7_else_1_else_acc_idiv[2:0];
  assign else_7_else_1_equal_tmp = g_1_lpi_dfm == mux1h_38_tmp;
  assign else_7_equal_tmp = r_1_lpi_dfm == mux1h_38_tmp;
  assign unequal_tmp_10 = (mux1h_38_tmp[9]) | (mux1h_38_tmp[8]) | (mux1h_38_tmp[7])
      | (mux1h_38_tmp[6]) | (mux1h_38_tmp[5]) | (mux1h_38_tmp[4]) | (mux1h_38_tmp[3])
      | (mux1h_38_tmp[2]) | (mux1h_38_tmp[1]) | (mux1h_38_tmp[0]);
  assign nl_if_3_acc_1_itm = ({1'b1 , g_rsc_mgc_in_wire_d , 1'b1}) + conv_u2u_11_12({(~
      r_rsc_mgc_in_wire_d) , 1'b1});
  assign if_3_acc_1_itm = nl_if_3_acc_1_itm[11:0];
  assign nl_if_acc_1_itm = ({1'b1 , r_rsc_mgc_in_wire_d , 1'b1}) + conv_u2u_11_12({(~
      g_rsc_mgc_in_wire_d) , 1'b1});
  assign if_acc_1_itm = nl_if_acc_1_itm[11:0];
  assign mux1h_40_nl = MUX1HOT_v_18_3_2({(div_mgc_div_16_z_oreg[17:0]) , (div_mgc_div_15_z_oreg[17:0])
      , s_sg1_1_sva_2_duc}, {(~((~(or_dcpl_807 | or_dcpl_805 | or_dcpl_803 | or_dcpl_801))
      | else_7_if_div_2cyc_st_3)) , ((or_dcpl_807 | or_dcpl_805 | or_dcpl_803 | or_dcpl_801)
      & else_7_if_div_2cyc_st_3) , ((~((max_sg1_lpi_dfm_3_st_3[9]) | (max_sg1_lpi_dfm_3_st_3[8])
      | (max_sg1_lpi_dfm_3_st_3[7]))) & (~((max_sg1_lpi_dfm_3_st_3[6]) | (max_sg1_lpi_dfm_3_st_3[5])))
      & (~((max_sg1_lpi_dfm_3_st_3[4]) | (max_sg1_lpi_dfm_3_st_3[3]) | (max_sg1_lpi_dfm_3_st_3[2])))
      & (~((max_sg1_lpi_dfm_3_st_3[1]) | (max_sg1_lpi_dfm_3_st_3[0]))))});
  assign nl_mul_1_itm = 18'b11001 * ((mux1h_40_nl) & ({{17{unequal_tmp_9}}, unequal_tmp_9})
      & ({{17{unequal_tmp_4}}, unequal_tmp_4}));
  assign mul_1_itm = nl_mul_1_itm[17:0];
  assign nl_mul_itm = 14'b11001 * conv_u2u_10_14(mux1h_38_tmp);
  assign mul_itm = nl_mul_itm[13:0];
  assign and_dcpl_23 = ~((else_7_if_1_div_5cyc_st_3[1]) | (else_7_if_1_div_5cyc_st_3[0]));
  assign and_dcpl_24 = main_stage_0_4 & else_7_equal_svs_st_3;
  assign and_dcpl_74 = ~((else_7_else_1_if_div_5cyc_st_3[2]) | (else_7_else_1_if_div_5cyc_st_3[1]));
  assign and_dcpl_76 = main_stage_0_4 & (~ else_7_equal_svs_st_3);
  assign and_dcpl_98 = (~ (else_7_else_1_if_div_5cyc_st_3[2])) & (else_7_else_1_if_div_5cyc_st_3[1]);
  assign and_dcpl_136 = ~((else_7_else_1_else_div_5cyc_st_3[1]) | (else_7_else_1_else_div_5cyc_st_3[2]));
  assign and_dcpl_160 = (else_7_else_1_else_div_5cyc_st_3[1]) & (~ (else_7_else_1_else_div_5cyc_st_3[2]));
  assign or_tmp_1 = (acc_2_psp_sva_st_2[0]) | (acc_2_psp_sva_st_2[9]) | (acc_2_psp_sva_st_2[8])
      | (acc_2_psp_sva_st_2[7]) | (acc_2_psp_sva_st_2[6]) | (acc_2_psp_sva_st_2[5])
      | (acc_2_psp_sva_st_2[4]) | (acc_2_psp_sva_st_2[3]) | (acc_2_psp_sva_st_2[2])
      | (acc_2_psp_sva_st_2[1]);
  assign and_dcpl_200 = ~((else_7_if_1_div_5cyc_st_2[1]) | (else_7_if_1_div_5cyc_st_2[0]));
  assign and_dcpl_201 = main_stage_0_3 & else_7_equal_svs_st_2;
  assign and_dcpl_241 = ~((else_7_else_1_if_div_5cyc_st_2[2]) | (else_7_else_1_if_div_5cyc_st_2[1]));
  assign and_dcpl_243 = main_stage_0_3 & (~ else_7_equal_svs_st_2);
  assign and_dcpl_261 = (~ (else_7_else_1_if_div_5cyc_st_2[2])) & (else_7_else_1_if_div_5cyc_st_2[1]);
  assign and_dcpl_293 = ~((else_7_else_1_else_div_5cyc_st_2[1]) | (else_7_else_1_else_div_5cyc_st_2[2]));
  assign and_dcpl_313 = (else_7_else_1_else_div_5cyc_st_2[1]) & (~ (else_7_else_1_else_div_5cyc_st_2[2]));
  assign and_dcpl_348 = main_stage_0_2 & else_7_equal_svs_st_1;
  assign and_dcpl_388 = ~((else_7_else_1_if_div_5cyc_st_1[2]) | (else_7_else_1_if_div_5cyc_st_1[1]));
  assign and_dcpl_408 = (~ (else_7_else_1_if_div_5cyc_st_1[2])) & (else_7_else_1_if_div_5cyc_st_1[1]);
  assign and_dcpl_440 = ~((else_7_else_1_else_div_5cyc_st_1[2]) | (else_7_else_1_else_div_5cyc_st_1[1]));
  assign and_dcpl_460 = (~ (else_7_else_1_else_div_5cyc_st_1[2])) & (else_7_else_1_else_div_5cyc_st_1[1]);
  assign or_tmp_3 = (else_7_if_1_acc_tmp[2]) | (else_7_if_1_acc_tmp[1]) | (else_7_if_1_acc_tmp[0]);
  assign or_tmp_11 = (else_7_if_1_acc_tmp[2]) | (else_7_if_1_acc_tmp[1]);
  assign or_tmp_79 = (else_7_else_1_else_acc_tmp[2]) | (else_7_else_1_else_acc_tmp[1])
      | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp | else_7_equal_tmp;
  assign and_dcpl_503 = ~((else_7_if_1_div_5cyc_st_5[0]) | (else_7_if_1_div_5cyc_st_5[2]));
  assign and_dcpl_504 = else_7_equal_svs_st_5 & (~ (else_7_if_1_div_5cyc_st_5[1]));
  assign and_dcpl_506 = (else_7_if_1_div_5cyc_st_5[0]) & (~ (else_7_if_1_div_5cyc_st_5[2]));
  assign and_dcpl_510 = else_7_equal_svs_st_5 & (else_7_if_1_div_5cyc_st_5[1]);
  assign and_dcpl_515 = (~ (else_7_if_1_div_5cyc_st_5[0])) & (else_7_if_1_div_5cyc_st_5[2]);
  assign and_dcpl_518 = ((else_7_if_1_div_5cyc_st_5[1]) | (else_7_if_1_div_5cyc_st_5[0]))
      & (else_7_if_1_div_5cyc_st_5[2]);
  assign and_dcpl_520 = main_stage_0_6 & else_7_equal_svs_st_5;
  assign and_dcpl_521 = and_dcpl_520 & (~ (else_7_if_1_div_5cyc_st_5[1]));
  assign and_dcpl_531 = and_dcpl_520 & (else_7_if_1_div_5cyc_st_5[1]);
  assign and_dcpl_554 = ~((else_7_else_1_if_div_5cyc_st_5[1]) | (else_7_else_1_if_div_5cyc_st_5[2]));
  assign and_dcpl_555 = (~ else_7_equal_svs_st_5) & else_7_else_1_equal_svs_st_5;
  assign and_dcpl_556 = and_dcpl_555 & (~ (else_7_else_1_if_div_5cyc_st_5[0]));
  assign and_dcpl_560 = and_dcpl_555 & (else_7_else_1_if_div_5cyc_st_5[0]);
  assign and_dcpl_562 = (else_7_else_1_if_div_5cyc_st_5[1]) & (~ (else_7_else_1_if_div_5cyc_st_5[2]));
  assign and_dcpl_574 = ((else_7_else_1_if_div_5cyc_st_5[0]) | (else_7_else_1_if_div_5cyc_st_5[1]))
      & (else_7_else_1_if_div_5cyc_st_5[2]);
  assign and_dcpl_575 = ~((else_7_else_1_if_div_5cyc_st_5[0]) | (else_7_else_1_if_div_5cyc_st_5[1]));
  assign and_588_cse = and_dcpl_575 & (~ (else_7_else_1_if_div_5cyc_st_5[2]));
  assign and_590_cse = (else_7_else_1_if_div_5cyc_st_5[0]) & (~ (else_7_else_1_if_div_5cyc_st_5[1]))
      & (~ (else_7_else_1_if_div_5cyc_st_5[2]));
  assign and_592_cse = (~ (else_7_else_1_if_div_5cyc_st_5[0])) & (else_7_else_1_if_div_5cyc_st_5[1])
      & (~ (else_7_else_1_if_div_5cyc_st_5[2]));
  assign and_594_cse = (else_7_else_1_if_div_5cyc_st_5[0]) & (else_7_else_1_if_div_5cyc_st_5[1])
      & (~ (else_7_else_1_if_div_5cyc_st_5[2]));
  assign and_596_cse = and_dcpl_575 & (else_7_else_1_if_div_5cyc_st_5[2]);
  assign and_dcpl_588 = main_stage_0_6 & (~ else_7_equal_svs_st_5);
  assign and_dcpl_589 = and_dcpl_588 & else_7_else_1_equal_svs_st_5;
  assign or_dcpl_462 = (~ main_stage_0_6) | else_7_equal_svs_st_5;
  assign and_dcpl_626 = ~((else_7_else_1_else_div_5cyc_st_5[0]) | (else_7_else_1_else_div_5cyc_st_5[2]));
  assign and_dcpl_627 = ~(else_7_equal_svs_st_5 | else_7_else_1_equal_svs_st_5);
  assign and_dcpl_628 = and_dcpl_627 & (~ (else_7_else_1_else_div_5cyc_st_5[1]));
  assign and_dcpl_630 = (else_7_else_1_else_div_5cyc_st_5[0]) & (~ (else_7_else_1_else_div_5cyc_st_5[2]));
  assign and_dcpl_636 = and_dcpl_627 & (else_7_else_1_else_div_5cyc_st_5[1]);
  assign and_dcpl_646 = ((else_7_else_1_else_div_5cyc_st_5[1]) | (else_7_else_1_else_div_5cyc_st_5[0]))
      & (else_7_else_1_else_div_5cyc_st_5[2]);
  assign and_dcpl_647 = ~((else_7_else_1_else_div_5cyc_st_5[1]) | (else_7_else_1_else_div_5cyc_st_5[0]));
  assign and_660_cse = and_dcpl_647 & (~ (else_7_else_1_else_div_5cyc_st_5[2]));
  assign and_662_cse = (~ (else_7_else_1_else_div_5cyc_st_5[1])) & (else_7_else_1_else_div_5cyc_st_5[0])
      & (~ (else_7_else_1_else_div_5cyc_st_5[2]));
  assign and_664_cse = (else_7_else_1_else_div_5cyc_st_5[1]) & (~ (else_7_else_1_else_div_5cyc_st_5[0]))
      & (~ (else_7_else_1_else_div_5cyc_st_5[2]));
  assign and_666_cse = (else_7_else_1_else_div_5cyc_st_5[1]) & (else_7_else_1_else_div_5cyc_st_5[0])
      & (~ (else_7_else_1_else_div_5cyc_st_5[2]));
  assign and_668_cse = and_dcpl_647 & (else_7_else_1_else_div_5cyc_st_5[2]);
  assign and_dcpl_661 = and_dcpl_588 & (~ else_7_else_1_equal_svs_st_5);
  assign and_dcpl_698 = ~((else_7_if_1_acc_tmp[1]) | (else_7_if_1_acc_tmp[0]));
  assign and_dcpl_699 = else_7_equal_tmp & (~ (else_7_if_1_acc_tmp[2]));
  assign and_dcpl_702 = ~((else_7_if_1_div_5cyc_st_1[0]) | (else_7_if_1_div_5cyc_st_1[1]));
  assign and_dcpl_704 = and_dcpl_348 & (~ (else_7_if_1_div_5cyc_st_1[2]));
  assign or_tmp_115 = (else_7_if_1_acc_tmp[0]) | (else_7_if_1_acc_tmp[1]) | (else_7_if_1_acc_tmp[2]);
  assign or_tmp_116 = (acc_2_psp_sva_st_1[1]) | (acc_2_psp_sva_st_1[2]) | (acc_2_psp_sva_st_1[3])
      | (acc_2_psp_sva_st_1[4]) | (acc_2_psp_sva_st_1[5]) | (acc_2_psp_sva_st_1[6])
      | (acc_2_psp_sva_st_1[7]) | (acc_2_psp_sva_st_1[8]) | (acc_2_psp_sva_st_1[9])
      | (acc_2_psp_sva_st_1[0]);
  assign nand_11_cse = ~(or_cse & else_7_equal_tmp);
  assign or_tmp_118 = ~(nand_11_cse & or_tmp_116);
  assign and_dcpl_709 = and_dcpl_201 & (~ (else_7_if_1_div_5cyc_st_2[2]));
  assign or_tmp_123 = ~((~(or_tmp_116 & main_stage_0_2)) & or_tmp_1);
  assign mux_236_nl = MUX_s_1_2_2({or_tmp_1 , (~ or_tmp_123)}, else_7_equal_svs_st_1);
  assign mux_tmp_35 = MUX_s_1_2_2({(mux_236_nl) , or_tmp_1}, (else_7_if_1_div_5cyc_st_1[1])
      | (else_7_if_1_div_5cyc_st_1[0]) | (else_7_if_1_div_5cyc_st_1[2]));
  assign and_dcpl_714 = and_dcpl_24 & (~ (else_7_if_1_div_5cyc_st_3[2]));
  assign or_tmp_126 = (acc_2_psp_sva_st_3[0]) | (acc_2_psp_sva_st_3[1]) | (acc_2_psp_sva_st_3[2])
      | (acc_2_psp_sva_st_3[3]) | (acc_2_psp_sva_st_3[4]) | (acc_2_psp_sva_st_3[5])
      | (acc_2_psp_sva_st_3[6]) | (acc_2_psp_sva_st_3[7]) | (acc_2_psp_sva_st_3[8])
      | (acc_2_psp_sva_st_3[9]);
  assign or_tmp_128 = (acc_2_psp_sva_st_1[0]) | (acc_2_psp_sva_st_1[1]) | (acc_2_psp_sva_st_1[2])
      | (acc_2_psp_sva_st_1[3]) | (acc_2_psp_sva_st_1[4]) | (acc_2_psp_sva_st_1[5])
      | (acc_2_psp_sva_st_1[6]) | (acc_2_psp_sva_st_1[7]) | (acc_2_psp_sva_st_1[8])
      | (acc_2_psp_sva_st_1[9]);
  assign or_tmp_130 = (acc_2_psp_sva_st_2[0]) | (acc_2_psp_sva_st_2[1]) | (acc_2_psp_sva_st_2[2])
      | (acc_2_psp_sva_st_2[3]) | (acc_2_psp_sva_st_2[4]) | (acc_2_psp_sva_st_2[5])
      | (acc_2_psp_sva_st_2[6]) | (acc_2_psp_sva_st_2[7]) | (acc_2_psp_sva_st_2[8])
      | (acc_2_psp_sva_st_2[9]);
  assign or_661_cse = (~ or_tmp_128) | (~ main_stage_0_2) | (~ else_7_equal_svs_st_1)
      | (else_7_if_1_div_5cyc_st_1[0]) | (else_7_if_1_div_5cyc_st_1[1]) | (else_7_if_1_div_5cyc_st_1[2]);
  assign or_663_cse = (~ or_tmp_130) | (~ main_stage_0_3) | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_5cyc_st_2[0]) | (else_7_if_1_div_5cyc_st_2[1]) | (else_7_if_1_div_5cyc_st_2[2]);
  assign and_tmp_1 = or_661_cse & or_663_cse;
  assign and_tmp_4 = or_661_cse & or_663_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | (~ else_7_equal_svs_st_3) | (else_7_if_1_div_5cyc_st_3[0]) | (else_7_if_1_div_5cyc_st_3[1])
      | (else_7_if_1_div_5cyc_st_3[2]));
  assign or_tmp_160 = (~ (else_7_if_1_acc_tmp[0])) | (else_7_if_1_acc_tmp[1]) | (else_7_if_1_acc_tmp[2]);
  assign mux_237_nl = MUX_s_1_2_2({or_tmp_1 , (~ or_tmp_123)}, else_7_equal_svs_st_1);
  assign mux_tmp_46 = MUX_s_1_2_2({(mux_237_nl) , or_tmp_1}, (else_7_if_1_div_5cyc_st_1[1])
      | (~ (else_7_if_1_div_5cyc_st_1[0])) | (else_7_if_1_div_5cyc_st_1[2]));
  assign or_718_cse = (~ or_tmp_128) | (~ main_stage_0_2) | (~ else_7_equal_svs_st_1)
      | (~ (else_7_if_1_div_5cyc_st_1[0])) | (else_7_if_1_div_5cyc_st_1[1]) | (else_7_if_1_div_5cyc_st_1[2]);
  assign or_720_cse = (~ or_tmp_130) | (~ main_stage_0_3) | (~ else_7_equal_svs_st_2)
      | (~ (else_7_if_1_div_5cyc_st_2[0])) | (else_7_if_1_div_5cyc_st_2[1]) | (else_7_if_1_div_5cyc_st_2[2]);
  assign and_tmp_9 = or_718_cse & or_720_cse;
  assign nor_tmp_10 = (else_7_if_1_acc_tmp[0]) & else_7_equal_tmp;
  assign and_tmp_12 = or_718_cse & or_720_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | (~ else_7_equal_svs_st_3) | (~ (else_7_if_1_div_5cyc_st_3[0])) | (else_7_if_1_div_5cyc_st_3[1])
      | (else_7_if_1_div_5cyc_st_3[2]));
  assign or_tmp_199 = (else_7_if_1_acc_tmp[0]) | (~ (else_7_if_1_acc_tmp[1])) | (else_7_if_1_acc_tmp[2]);
  assign mux_238_nl = MUX_s_1_2_2({or_tmp_1 , (~ or_tmp_123)}, else_7_equal_svs_st_1);
  assign mux_tmp_57 = MUX_s_1_2_2({(mux_238_nl) , or_tmp_1}, (~ (else_7_if_1_div_5cyc_st_1[1]))
      | (else_7_if_1_div_5cyc_st_1[0]) | (else_7_if_1_div_5cyc_st_1[2]));
  assign or_tmp_205 = (else_7_if_1_acc_tmp[2]) | (~ (else_7_if_1_acc_tmp[1])) | (else_7_if_1_acc_tmp[0]);
  assign or_775_cse = (~ or_tmp_128) | (~ main_stage_0_2) | (~ else_7_equal_svs_st_1)
      | (else_7_if_1_div_5cyc_st_1[0]) | (~ (else_7_if_1_div_5cyc_st_1[1])) | (else_7_if_1_div_5cyc_st_1[2]);
  assign or_777_cse = (~ or_tmp_130) | (~ main_stage_0_3) | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_5cyc_st_2[0]) | (~ (else_7_if_1_div_5cyc_st_2[1])) | (else_7_if_1_div_5cyc_st_2[2]);
  assign and_tmp_17 = or_775_cse & or_777_cse;
  assign and_tmp_20 = or_775_cse & or_777_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | (~ else_7_equal_svs_st_3) | (else_7_if_1_div_5cyc_st_3[0]) | (~ (else_7_if_1_div_5cyc_st_3[1]))
      | (else_7_if_1_div_5cyc_st_3[2]));
  assign or_tmp_238 = (~ (else_7_if_1_acc_tmp[0])) | (~ (else_7_if_1_acc_tmp[1]))
      | (else_7_if_1_acc_tmp[2]);
  assign mux_89_nl = MUX_s_1_2_2({or_tmp_1 , (~ or_tmp_123)}, else_7_equal_svs_st_1);
  assign mux_tmp_68 = MUX_s_1_2_2({(mux_89_nl) , or_tmp_1}, (~ (else_7_if_1_div_5cyc_st_1[1]))
      | (~ (else_7_if_1_div_5cyc_st_1[0])) | (else_7_if_1_div_5cyc_st_1[2]));
  assign nand_22_cse = ~(or_tmp_128 & main_stage_0_2 & else_7_equal_svs_st_1 & (else_7_if_1_div_5cyc_st_1[0])
      & (else_7_if_1_div_5cyc_st_1[1]) & (~ (else_7_if_1_div_5cyc_st_1[2])));
  assign nand_23_cse = ~(or_tmp_130 & main_stage_0_3 & else_7_equal_svs_st_2 & (else_7_if_1_div_5cyc_st_2[0])
      & (else_7_if_1_div_5cyc_st_2[1]) & (~ (else_7_if_1_div_5cyc_st_2[2])));
  assign and_tmp_25 = nand_22_cse & nand_23_cse;
  assign nor_tmp_16 = (else_7_if_1_acc_tmp[1]) & (else_7_if_1_acc_tmp[0]) & else_7_equal_tmp;
  assign and_tmp_28 = nand_22_cse & nand_23_cse & (~(or_tmp_126 & main_stage_0_4
      & else_7_equal_svs_st_3 & (else_7_if_1_div_5cyc_st_3[0]) & (else_7_if_1_div_5cyc_st_3[1])
      & (~ (else_7_if_1_div_5cyc_st_3[2]))));
  assign or_tmp_273 = (else_7_if_1_acc_tmp[0]) | (else_7_if_1_acc_tmp[1]);
  assign mux_135_nl = MUX_s_1_2_2({or_tmp_1 , (~ or_tmp_123)}, (else_7_if_1_div_5cyc_st_1[2])
      & else_7_equal_svs_st_1);
  assign mux_tmp_81 = MUX_s_1_2_2({(mux_135_nl) , or_tmp_1}, (else_7_if_1_div_5cyc_st_1[1])
      | (else_7_if_1_div_5cyc_st_1[0]));
  assign or_tmp_279 = (~ (else_7_if_1_acc_tmp[2])) | (else_7_if_1_acc_tmp[1]) | (else_7_if_1_acc_tmp[0]);
  assign or_tmp_284 = (~ or_tmp_130) | (~ main_stage_0_3) | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_5cyc_st_2[0]) | (else_7_if_1_div_5cyc_st_2[1]) | (~ (else_7_if_1_div_5cyc_st_2[2]));
  assign or_885_cse = (~ or_tmp_128) | (~ main_stage_0_2) | (~ else_7_equal_svs_st_1)
      | (else_7_if_1_div_5cyc_st_1[0]) | (else_7_if_1_div_5cyc_st_1[1]);
  assign mux_tmp_84 = MUX_s_1_2_2({(~((else_7_if_1_div_5cyc_st_1[2]) | (~ or_tmp_284)))
      , or_tmp_284}, or_885_cse);
  assign or_tmp_295 = (~ or_tmp_126) | (~ main_stage_0_4) | (~ else_7_equal_svs_st_3)
      | (else_7_if_1_div_5cyc_st_3[0]) | (else_7_if_1_div_5cyc_st_3[1]) | (~ (else_7_if_1_div_5cyc_st_3[2]));
  assign mux_tmp_87 = MUX_s_1_2_2({(~((else_7_if_1_div_5cyc_st_2[2]) | (~ or_tmp_295)))
      , or_tmp_295}, (~ or_tmp_130) | (~ main_stage_0_3) | (~ else_7_equal_svs_st_2)
      | (else_7_if_1_div_5cyc_st_2[0]) | (else_7_if_1_div_5cyc_st_2[1]));
  assign mux_143_cse = MUX_s_1_2_2({(~((else_7_if_1_div_5cyc_st_1[2]) | (~ mux_tmp_87)))
      , mux_tmp_87}, or_885_cse);
  assign and_dcpl_888 = ~((else_7_else_1_if_acc_tmp[1]) | (else_7_else_1_if_acc_tmp[0]));
  assign and_dcpl_889 = (~ else_7_equal_tmp) & else_7_else_1_equal_tmp;
  assign and_dcpl_890 = and_dcpl_889 & (~ (else_7_else_1_if_acc_tmp[2]));
  assign and_dcpl_896 = and_504_cse & else_7_else_1_equal_svs_st_1;
  assign or_tmp_322 = (else_7_else_1_if_acc_tmp[0]) | (else_7_else_1_if_acc_tmp[1])
      | (else_7_else_1_if_acc_tmp[2]);
  assign or_946_cse = (~ or_cse) | (~ else_7_else_1_equal_tmp) | else_7_equal_tmp;
  assign and_tmp_35 = or_946_cse & or_tmp_116;
  assign mux_tmp_99 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (else_7_else_1_if_div_5cyc_st_1[0])
      | (else_7_else_1_if_div_5cyc_st_1[1]) | (else_7_else_1_if_div_5cyc_st_1[2])
      | (~ else_7_else_1_equal_svs_st_1) | else_7_equal_svs_st_1);
  assign or_tmp_330 = (else_7_else_1_if_acc_tmp[2]) | (else_7_else_1_if_acc_tmp[1])
      | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp) | else_7_equal_tmp;
  assign or_954_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | (~ else_7_else_1_equal_svs_st_1) | (else_7_else_1_if_div_5cyc_st_1[0]) |
      (else_7_else_1_if_div_5cyc_st_1[1]) | (else_7_else_1_if_div_5cyc_st_1[2]);
  assign or_956_cse = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_5cyc_st_2[0]) |
      (else_7_else_1_if_div_5cyc_st_2[1]) | (else_7_else_1_if_div_5cyc_st_2[2]);
  assign and_tmp_37 = or_954_cse & or_956_cse;
  assign and_tmp_40 = or_954_cse & or_956_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | else_7_equal_svs_st_3 | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_5cyc_st_3[0])
      | (else_7_else_1_if_div_5cyc_st_3[1]) | (else_7_else_1_if_div_5cyc_st_3[2]));
  assign or_tmp_363 = (~ (else_7_else_1_if_acc_tmp[0])) | (else_7_else_1_if_acc_tmp[1])
      | (else_7_else_1_if_acc_tmp[2]);
  assign mux_tmp_106 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (~ (else_7_else_1_if_div_5cyc_st_1[0]))
      | (else_7_else_1_if_div_5cyc_st_1[1]) | (else_7_else_1_if_div_5cyc_st_1[2])
      | (~ else_7_else_1_equal_svs_st_1) | else_7_equal_svs_st_1);
  assign or_tmp_369 = (else_7_else_1_if_acc_tmp[2]) | (else_7_else_1_if_acc_tmp[1])
      | (~ (else_7_else_1_if_acc_tmp[0])) | (~ else_7_else_1_equal_tmp) | else_7_equal_tmp;
  assign or_1011_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | (~ else_7_else_1_equal_svs_st_1) | (~ (else_7_else_1_if_div_5cyc_st_1[0]))
      | (else_7_else_1_if_div_5cyc_st_1[1]) | (else_7_else_1_if_div_5cyc_st_1[2]);
  assign or_1013_cse = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (~ (else_7_else_1_if_div_5cyc_st_2[0]))
      | (else_7_else_1_if_div_5cyc_st_2[1]) | (else_7_else_1_if_div_5cyc_st_2[2]);
  assign and_tmp_46 = or_1011_cse & or_1013_cse;
  assign and_tmp_49 = or_1011_cse & or_1013_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | else_7_equal_svs_st_3 | (~ else_7_else_1_equal_svs_st_3) | (~ (else_7_else_1_if_div_5cyc_st_3[0]))
      | (else_7_else_1_if_div_5cyc_st_3[1]) | (else_7_else_1_if_div_5cyc_st_3[2]));
  assign or_tmp_402 = (else_7_else_1_if_acc_tmp[0]) | (~ (else_7_else_1_if_acc_tmp[1]))
      | (else_7_else_1_if_acc_tmp[2]);
  assign mux_tmp_113 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (else_7_else_1_if_div_5cyc_st_1[0])
      | (~ (else_7_else_1_if_div_5cyc_st_1[1])) | (else_7_else_1_if_div_5cyc_st_1[2])
      | (~ else_7_else_1_equal_svs_st_1) | else_7_equal_svs_st_1);
  assign or_tmp_408 = (else_7_else_1_if_acc_tmp[2]) | (~ (else_7_else_1_if_acc_tmp[1]))
      | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp) | else_7_equal_tmp;
  assign or_1068_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | (~ else_7_else_1_equal_svs_st_1) | (else_7_else_1_if_div_5cyc_st_1[0]) |
      (~ (else_7_else_1_if_div_5cyc_st_1[1])) | (else_7_else_1_if_div_5cyc_st_1[2]);
  assign or_1070_cse = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_5cyc_st_2[0]) |
      (~ (else_7_else_1_if_div_5cyc_st_2[1])) | (else_7_else_1_if_div_5cyc_st_2[2]);
  assign and_tmp_55 = or_1068_cse & or_1070_cse;
  assign and_tmp_58 = or_1068_cse & or_1070_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | else_7_equal_svs_st_3 | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_5cyc_st_3[0])
      | (~ (else_7_else_1_if_div_5cyc_st_3[1])) | (else_7_else_1_if_div_5cyc_st_3[2]));
  assign or_tmp_441 = (~ (else_7_else_1_if_acc_tmp[0])) | (~ (else_7_else_1_if_acc_tmp[1]))
      | (else_7_else_1_if_acc_tmp[2]);
  assign mux_tmp_120 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (~ (else_7_else_1_if_div_5cyc_st_1[0]))
      | (~ (else_7_else_1_if_div_5cyc_st_1[1])) | (else_7_else_1_if_div_5cyc_st_1[2])
      | (~ else_7_else_1_equal_svs_st_1) | else_7_equal_svs_st_1);
  assign or_tmp_447 = (else_7_else_1_if_acc_tmp[2]) | (~ (else_7_else_1_if_acc_tmp[1]))
      | (~ (else_7_else_1_if_acc_tmp[0])) | (~ else_7_else_1_equal_tmp) | else_7_equal_tmp;
  assign nand_34_cse = ~(or_tmp_128 & main_stage_0_2 & (~ else_7_equal_svs_st_1)
      & else_7_else_1_equal_svs_st_1 & (else_7_else_1_if_div_5cyc_st_1[0]) & (else_7_else_1_if_div_5cyc_st_1[1])
      & (~ (else_7_else_1_if_div_5cyc_st_1[2])));
  assign nand_35_cse = ~(or_tmp_130 & main_stage_0_3 & (~ else_7_equal_svs_st_2)
      & else_7_else_1_equal_svs_st_2 & (else_7_else_1_if_div_5cyc_st_2[0]) & (else_7_else_1_if_div_5cyc_st_2[1])
      & (~ (else_7_else_1_if_div_5cyc_st_2[2])));
  assign and_tmp_64 = nand_34_cse & nand_35_cse;
  assign and_tmp_67 = nand_34_cse & nand_35_cse & (~(or_tmp_126 & main_stage_0_4
      & (~ else_7_equal_svs_st_3) & else_7_else_1_equal_svs_st_3 & (else_7_else_1_if_div_5cyc_st_3[0])
      & (else_7_else_1_if_div_5cyc_st_3[1]) & (~ (else_7_else_1_if_div_5cyc_st_3[2]))));
  assign nor_tmp_22 = ~((else_7_else_1_if_acc_tmp[0]) | (else_7_else_1_if_acc_tmp[1])
      | (~ (else_7_else_1_if_acc_tmp[2])));
  assign mux_tmp_127 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (else_7_else_1_if_div_5cyc_st_1[0])
      | (else_7_else_1_if_div_5cyc_st_1[1]) | (~ (else_7_else_1_if_div_5cyc_st_1[2]))
      | (~ else_7_else_1_equal_svs_st_1) | else_7_equal_svs_st_1);
  assign or_tmp_484 = (~ (else_7_else_1_if_acc_tmp[2])) | (else_7_else_1_if_acc_tmp[1])
      | (else_7_else_1_if_acc_tmp[0]) | (~ else_7_else_1_equal_tmp) | else_7_equal_tmp;
  assign or_tmp_489 = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_5cyc_st_2[0]) |
      (else_7_else_1_if_div_5cyc_st_2[1]) | (~ (else_7_else_1_if_div_5cyc_st_2[2]));
  assign or_1180_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | (~ else_7_else_1_equal_svs_st_1) | (else_7_else_1_if_div_5cyc_st_1[0]) |
      (else_7_else_1_if_div_5cyc_st_1[1]);
  assign mux_tmp_129 = MUX_s_1_2_2({(~((else_7_else_1_if_div_5cyc_st_1[2]) | (~ or_tmp_489)))
      , or_tmp_489}, or_1180_cse);
  assign or_tmp_500 = (~ or_tmp_126) | (~ main_stage_0_4) | else_7_equal_svs_st_3
      | (~ else_7_else_1_equal_svs_st_3) | (else_7_else_1_if_div_5cyc_st_3[0]) |
      (else_7_else_1_if_div_5cyc_st_3[1]) | (~ (else_7_else_1_if_div_5cyc_st_3[2]));
  assign mux_tmp_131 = MUX_s_1_2_2({(~((else_7_else_1_if_div_5cyc_st_2[2]) | (~ or_tmp_500)))
      , or_tmp_500}, (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | (~ else_7_else_1_equal_svs_st_2) | (else_7_else_1_if_div_5cyc_st_2[0]) |
      (else_7_else_1_if_div_5cyc_st_2[1]));
  assign mux_187_cse = MUX_s_1_2_2({(~((else_7_else_1_if_div_5cyc_st_1[2]) | (~ mux_tmp_131)))
      , mux_tmp_131}, or_1180_cse);
  assign and_dcpl_1118 = ~((else_7_else_1_else_acc_tmp[1]) | (else_7_else_1_else_acc_tmp[0]));
  assign and_dcpl_1119 = ~(else_7_equal_tmp | else_7_else_1_equal_tmp);
  assign and_dcpl_1120 = and_dcpl_1119 & (~ (else_7_else_1_else_acc_tmp[2]));
  assign and_dcpl_1126 = and_504_cse & (~ else_7_else_1_equal_svs_st_1);
  assign or_tmp_527 = (else_7_else_1_else_acc_tmp[0]) | (else_7_else_1_else_acc_tmp[1])
      | (else_7_else_1_else_acc_tmp[2]);
  assign or_1241_cse = (~ or_cse) | else_7_else_1_equal_tmp | else_7_equal_tmp;
  assign and_tmp_75 = or_1241_cse & or_tmp_116;
  assign mux_tmp_140 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (else_7_else_1_else_div_5cyc_st_1[0])
      | (else_7_else_1_else_div_5cyc_st_1[1]) | (else_7_else_1_else_div_5cyc_st_1[2])
      | else_7_else_1_equal_svs_st_1 | else_7_equal_svs_st_1);
  assign or_1249_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | else_7_else_1_equal_svs_st_1 | (else_7_else_1_else_div_5cyc_st_1[0]) | (else_7_else_1_else_div_5cyc_st_1[1])
      | (else_7_else_1_else_div_5cyc_st_1[2]);
  assign or_1251_cse = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_5cyc_st_2[0]) | (else_7_else_1_else_div_5cyc_st_2[1])
      | (else_7_else_1_else_div_5cyc_st_2[2]);
  assign and_tmp_77 = or_1249_cse & or_1251_cse;
  assign and_tmp_80 = or_1249_cse & or_1251_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | else_7_equal_svs_st_3 | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_5cyc_st_3[0])
      | (else_7_else_1_else_div_5cyc_st_3[1]) | (else_7_else_1_else_div_5cyc_st_3[2]));
  assign or_tmp_568 = (~ (else_7_else_1_else_acc_tmp[0])) | (else_7_else_1_else_acc_tmp[1])
      | (else_7_else_1_else_acc_tmp[2]);
  assign mux_tmp_147 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (~ (else_7_else_1_else_div_5cyc_st_1[0]))
      | (else_7_else_1_else_div_5cyc_st_1[1]) | (else_7_else_1_else_div_5cyc_st_1[2])
      | else_7_else_1_equal_svs_st_1 | else_7_equal_svs_st_1);
  assign or_tmp_574 = (else_7_else_1_else_acc_tmp[2]) | (else_7_else_1_else_acc_tmp[1])
      | (~ (else_7_else_1_else_acc_tmp[0])) | else_7_else_1_equal_tmp | else_7_equal_tmp;
  assign or_1306_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | else_7_else_1_equal_svs_st_1 | (~ (else_7_else_1_else_div_5cyc_st_1[0]))
      | (else_7_else_1_else_div_5cyc_st_1[1]) | (else_7_else_1_else_div_5cyc_st_1[2]);
  assign or_1308_cse = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (~ (else_7_else_1_else_div_5cyc_st_2[0]))
      | (else_7_else_1_else_div_5cyc_st_2[1]) | (else_7_else_1_else_div_5cyc_st_2[2]);
  assign and_tmp_86 = or_1306_cse & or_1308_cse;
  assign and_tmp_89 = or_1306_cse & or_1308_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | else_7_equal_svs_st_3 | else_7_else_1_equal_svs_st_3 | (~ (else_7_else_1_else_div_5cyc_st_3[0]))
      | (else_7_else_1_else_div_5cyc_st_3[1]) | (else_7_else_1_else_div_5cyc_st_3[2]));
  assign or_tmp_607 = (else_7_else_1_else_acc_tmp[0]) | (~ (else_7_else_1_else_acc_tmp[1]))
      | (else_7_else_1_else_acc_tmp[2]);
  assign mux_tmp_154 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (else_7_else_1_else_div_5cyc_st_1[0])
      | (~ (else_7_else_1_else_div_5cyc_st_1[1])) | (else_7_else_1_else_div_5cyc_st_1[2])
      | else_7_else_1_equal_svs_st_1 | else_7_equal_svs_st_1);
  assign or_tmp_613 = (else_7_else_1_else_acc_tmp[2]) | (~ (else_7_else_1_else_acc_tmp[1]))
      | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp | else_7_equal_tmp;
  assign or_1363_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | else_7_else_1_equal_svs_st_1 | (else_7_else_1_else_div_5cyc_st_1[0]) | (~
      (else_7_else_1_else_div_5cyc_st_1[1])) | (else_7_else_1_else_div_5cyc_st_1[2]);
  assign or_1365_cse = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_5cyc_st_2[0]) | (~
      (else_7_else_1_else_div_5cyc_st_2[1])) | (else_7_else_1_else_div_5cyc_st_2[2]);
  assign and_tmp_95 = or_1363_cse & or_1365_cse;
  assign and_tmp_98 = or_1363_cse & or_1365_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | else_7_equal_svs_st_3 | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_5cyc_st_3[0])
      | (~ (else_7_else_1_else_div_5cyc_st_3[1])) | (else_7_else_1_else_div_5cyc_st_3[2]));
  assign or_tmp_646 = (~ (else_7_else_1_else_acc_tmp[0])) | (~ (else_7_else_1_else_acc_tmp[1]))
      | (else_7_else_1_else_acc_tmp[2]);
  assign mux_tmp_161 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (~ (else_7_else_1_else_div_5cyc_st_1[0]))
      | (~ (else_7_else_1_else_div_5cyc_st_1[1])) | (else_7_else_1_else_div_5cyc_st_1[2])
      | else_7_else_1_equal_svs_st_1 | else_7_equal_svs_st_1);
  assign or_tmp_652 = (else_7_else_1_else_acc_tmp[2]) | (~ (else_7_else_1_else_acc_tmp[1]))
      | (~ (else_7_else_1_else_acc_tmp[0])) | else_7_else_1_equal_tmp | else_7_equal_tmp;
  assign or_1420_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | else_7_else_1_equal_svs_st_1 | (~ (else_7_else_1_else_div_5cyc_st_1[0]))
      | (~ (else_7_else_1_else_div_5cyc_st_1[1])) | (else_7_else_1_else_div_5cyc_st_1[2]);
  assign or_1422_cse = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (~ (else_7_else_1_else_div_5cyc_st_2[0]))
      | (~ (else_7_else_1_else_div_5cyc_st_2[1])) | (else_7_else_1_else_div_5cyc_st_2[2]);
  assign and_tmp_104 = or_1420_cse & or_1422_cse;
  assign and_tmp_107 = or_1420_cse & or_1422_cse & ((~ or_tmp_126) | (~ main_stage_0_4)
      | else_7_equal_svs_st_3 | else_7_else_1_equal_svs_st_3 | (~ (else_7_else_1_else_div_5cyc_st_3[0]))
      | (~ (else_7_else_1_else_div_5cyc_st_3[1])) | (else_7_else_1_else_div_5cyc_st_3[2]));
  assign nor_tmp_24 = ~((else_7_else_1_else_acc_tmp[0]) | (else_7_else_1_else_acc_tmp[1])
      | (~ (else_7_else_1_else_acc_tmp[2])));
  assign mux_tmp_168 = MUX_s_1_2_2({(~ or_tmp_123) , or_tmp_1}, (else_7_else_1_else_div_5cyc_st_1[0])
      | (else_7_else_1_else_div_5cyc_st_1[1]) | (~ (else_7_else_1_else_div_5cyc_st_1[2]))
      | else_7_else_1_equal_svs_st_1 | else_7_equal_svs_st_1);
  assign or_tmp_689 = (~ (else_7_else_1_else_acc_tmp[2])) | (else_7_else_1_else_acc_tmp[1])
      | (else_7_else_1_else_acc_tmp[0]) | else_7_else_1_equal_tmp | else_7_equal_tmp;
  assign or_tmp_694 = (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_5cyc_st_2[0]) | (else_7_else_1_else_div_5cyc_st_2[1])
      | (~ (else_7_else_1_else_div_5cyc_st_2[2]));
  assign or_1475_cse = (~ or_tmp_128) | (~ main_stage_0_2) | else_7_equal_svs_st_1
      | else_7_else_1_equal_svs_st_1 | (else_7_else_1_else_div_5cyc_st_1[0]) | (else_7_else_1_else_div_5cyc_st_1[1]);
  assign mux_tmp_170 = MUX_s_1_2_2({(~((else_7_else_1_else_div_5cyc_st_1[2]) | (~
      or_tmp_694))) , or_tmp_694}, or_1475_cse);
  assign or_tmp_705 = (~ or_tmp_126) | (~ main_stage_0_4) | else_7_equal_svs_st_3
      | else_7_else_1_equal_svs_st_3 | (else_7_else_1_else_div_5cyc_st_3[0]) | (else_7_else_1_else_div_5cyc_st_3[1])
      | (~ (else_7_else_1_else_div_5cyc_st_3[2]));
  assign mux_tmp_172 = MUX_s_1_2_2({(~((else_7_else_1_else_div_5cyc_st_2[2]) | (~
      or_tmp_705))) , or_tmp_705}, (~ or_tmp_130) | (~ main_stage_0_3) | else_7_equal_svs_st_2
      | else_7_else_1_equal_svs_st_2 | (else_7_else_1_else_div_5cyc_st_2[0]) | (else_7_else_1_else_div_5cyc_st_2[1]));
  assign mux_228_cse = MUX_s_1_2_2({(~((else_7_else_1_else_div_5cyc_st_1[2]) | (~
      mux_tmp_172))) , mux_tmp_172}, or_1475_cse);
  assign not_tmp_349 = ~(((mux1h_38_tmp[9]) | (mux1h_38_tmp[8]) | (mux1h_38_tmp[7])
      | (mux1h_38_tmp[6]) | (mux1h_38_tmp[5]) | (mux1h_38_tmp[4]) | (mux1h_38_tmp[3])
      | (mux1h_38_tmp[2]) | (mux1h_38_tmp[1]) | (mux1h_38_tmp[0])) & or_cse);
  assign or_dcpl_790 = not_tmp_349 | (~ else_7_if_div_2cyc);
  assign or_dcpl_792 = not_tmp_349 | else_7_if_div_2cyc;
  assign and_dcpl_1348 = ~((acc_itm[9]) | (acc_itm[10]));
  assign and_dcpl_1350 = ~((acc_itm[6]) | (acc_itm[7]) | (acc_itm[8]));
  assign and_dcpl_1352 = ~((acc_itm[4]) | (acc_itm[5]));
  assign and_dcpl_1354 = ~((acc_itm[1]) | (acc_itm[2]) | (acc_itm[3]));
  assign or_dcpl_801 = (max_sg1_lpi_dfm_3_st_3[1]) | (max_sg1_lpi_dfm_3_st_3[0]);
  assign or_dcpl_803 = (max_sg1_lpi_dfm_3_st_3[4]) | (max_sg1_lpi_dfm_3_st_3[3])
      | (max_sg1_lpi_dfm_3_st_3[2]);
  assign or_dcpl_805 = (max_sg1_lpi_dfm_3_st_3[6]) | (max_sg1_lpi_dfm_3_st_3[5]);
  assign or_dcpl_807 = (max_sg1_lpi_dfm_3_st_3[9]) | (max_sg1_lpi_dfm_3_st_3[8])
      | (max_sg1_lpi_dfm_3_st_3[7]);
  assign and_tmp_116 = ((max_sg1_lpi_dfm_3_st_3[0]) | (max_sg1_lpi_dfm_3_st_3[1])
      | (max_sg1_lpi_dfm_3_st_3[2]) | (max_sg1_lpi_dfm_3_st_3[3]) | (max_sg1_lpi_dfm_3_st_3[4])
      | (max_sg1_lpi_dfm_3_st_3[5]) | (max_sg1_lpi_dfm_3_st_3[6]) | (max_sg1_lpi_dfm_3_st_3[7])
      | (max_sg1_lpi_dfm_3_st_3[8]) | (max_sg1_lpi_dfm_3_st_3[9])) & ((acc_2_psp_sva_st_3[1])
      | (acc_2_psp_sva_st_3[9]) | (acc_2_psp_sva_st_3[8]) | (acc_2_psp_sva_st_3[7])
      | (acc_2_psp_sva_st_3[6]) | (acc_2_psp_sva_st_3[5]) | (acc_2_psp_sva_st_3[4])
      | (acc_2_psp_sva_st_3[3]) | (acc_2_psp_sva_st_3[2]) | (acc_2_psp_sva_st_3[0]));
  assign mux_92_nl = MUX_s_1_2_2({and_tmp_1 , (~(or_cse | (~ and_tmp_1)))}, else_7_equal_tmp);
  assign mux_93_nl = MUX_s_1_2_2({(mux_92_nl) , and_tmp_1}, or_tmp_3);
  assign and_730_cse = or_tmp_126 & (mux_93_nl) & and_dcpl_714 & and_dcpl_23;
  assign mux_94_nl = MUX_s_1_2_2({and_tmp_4 , (~(or_cse | (~ and_tmp_4)))}, else_7_equal_tmp);
  assign mux_95_cse = MUX_s_1_2_2({(mux_94_nl) , and_tmp_4}, or_tmp_3);
  assign mux_103_nl = MUX_s_1_2_2({and_tmp_9 , (~(or_cse | (~ and_tmp_9)))}, nor_tmp_10);
  assign mux_104_nl = MUX_s_1_2_2({(mux_103_nl) , and_tmp_9}, or_tmp_11);
  assign and_776_cse = or_tmp_126 & (mux_104_nl) & and_dcpl_714 & (~ (else_7_if_1_div_5cyc_st_3[1]))
      & (else_7_if_1_div_5cyc_st_3[0]);
  assign mux_105_nl = MUX_s_1_2_2({and_tmp_12 , (~(or_cse | (~ and_tmp_12)))}, nor_tmp_10);
  assign mux_106_cse = MUX_s_1_2_2({(mux_105_nl) , and_tmp_12}, or_tmp_11);
  assign mux_114_nl = MUX_s_1_2_2({and_tmp_17 , (~(or_cse | (~ and_tmp_17)))}, else_7_equal_tmp);
  assign mux_115_nl = MUX_s_1_2_2({(mux_114_nl) , and_tmp_17}, or_tmp_205);
  assign and_822_cse = or_tmp_126 & (mux_115_nl) & and_dcpl_714 & (else_7_if_1_div_5cyc_st_3[1])
      & (~ (else_7_if_1_div_5cyc_st_3[0]));
  assign mux_116_nl = MUX_s_1_2_2({and_tmp_20 , (~(or_cse | (~ and_tmp_20)))}, else_7_equal_tmp);
  assign mux_117_cse = MUX_s_1_2_2({(mux_116_nl) , and_tmp_20}, or_tmp_205);
  assign mux_125_nl = MUX_s_1_2_2({and_tmp_25 , (~(or_cse | (~ and_tmp_25)))}, nor_tmp_16);
  assign mux_126_nl = MUX_s_1_2_2({(mux_125_nl) , and_tmp_25}, else_7_if_1_acc_tmp[2]);
  assign and_868_cse = or_tmp_126 & (mux_126_nl) & and_dcpl_714 & (else_7_if_1_div_5cyc_st_3[1])
      & (else_7_if_1_div_5cyc_st_3[0]);
  assign mux_127_nl = MUX_s_1_2_2({and_tmp_28 , (~(or_cse | (~ and_tmp_28)))}, nor_tmp_16);
  assign mux_128_cse = MUX_s_1_2_2({(mux_127_nl) , and_tmp_28}, else_7_if_1_acc_tmp[2]);
  assign mux_140_nl = MUX_s_1_2_2({mux_tmp_84 , (~(or_cse | (~ mux_tmp_84)))}, else_7_equal_tmp);
  assign mux_141_nl = MUX_s_1_2_2({(mux_140_nl) , mux_tmp_84}, or_tmp_279);
  assign and_913_cse = or_tmp_126 & (mux_141_nl) & and_dcpl_24 & (else_7_if_1_div_5cyc_st_3[2])
      & and_dcpl_23;
  assign mux_144_nl = MUX_s_1_2_2({mux_143_cse , (~(or_cse | (~ mux_143_cse)))},
      else_7_equal_tmp);
  assign mux_145_cse = MUX_s_1_2_2({(mux_144_nl) , mux_143_cse}, or_tmp_279);
  assign mux_156_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_37))) , and_tmp_37}, or_tmp_330);
  assign and_960_cse = or_tmp_126 & (mux_156_nl) & and_146_cse & and_dcpl_74 & (~
      (else_7_else_1_if_div_5cyc_st_3[0]));
  assign mux_157_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_40))) , and_tmp_40}, or_tmp_330);
  assign mux_163_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_46))) , and_tmp_46}, or_tmp_369);
  assign and_1015_cse = or_tmp_126 & (mux_163_nl) & and_146_cse & and_dcpl_74 & (else_7_else_1_if_div_5cyc_st_3[0]);
  assign mux_164_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_49))) , and_tmp_49}, or_tmp_369);
  assign mux_170_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_55))) , and_tmp_55}, or_tmp_408);
  assign and_1070_cse = or_tmp_126 & (mux_170_nl) & and_146_cse & and_dcpl_98 & (~
      (else_7_else_1_if_div_5cyc_st_3[0]));
  assign mux_171_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_58))) , and_tmp_58}, or_tmp_408);
  assign mux_177_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_64))) , and_tmp_64}, or_tmp_447);
  assign and_1125_cse = or_tmp_126 & (mux_177_nl) & and_146_cse & and_dcpl_98 & (else_7_else_1_if_div_5cyc_st_3[0]);
  assign mux_178_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_67))) , and_tmp_67}, or_tmp_447);
  assign mux_185_nl = MUX_s_1_2_2({(~(or_cse | (~ mux_tmp_129))) , mux_tmp_129},
      or_tmp_484);
  assign and_1179_cse = or_tmp_126 & (mux_185_nl) & and_146_cse & (else_7_else_1_if_div_5cyc_st_3[2])
      & (~ (else_7_else_1_if_div_5cyc_st_3[1])) & (~ (else_7_else_1_if_div_5cyc_st_3[0]));
  assign mux_188_cse = MUX_s_1_2_2({(~(or_cse | (~ mux_187_cse))) , mux_187_cse},
      or_tmp_484);
  assign mux_197_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_77))) , and_tmp_77}, or_tmp_79);
  assign and_1230_cse = or_tmp_126 & (mux_197_nl) & and_208_cse & and_dcpl_136 &
      (~ (else_7_else_1_else_div_5cyc_st_3[0]));
  assign mux_198_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_80))) , and_tmp_80}, or_tmp_79);
  assign mux_204_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_86))) , and_tmp_86}, or_tmp_574);
  assign and_1285_cse = or_tmp_126 & (mux_204_nl) & and_208_cse & and_dcpl_136 &
      (else_7_else_1_else_div_5cyc_st_3[0]);
  assign mux_205_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_89))) , and_tmp_89}, or_tmp_574);
  assign mux_211_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_95))) , and_tmp_95}, or_tmp_613);
  assign and_1340_cse = or_tmp_126 & (mux_211_nl) & and_208_cse & and_dcpl_160 &
      (~ (else_7_else_1_else_div_5cyc_st_3[0]));
  assign mux_212_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_98))) , and_tmp_98}, or_tmp_613);
  assign mux_218_nl = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_104))) , and_tmp_104},
      or_tmp_652);
  assign and_1395_cse = or_tmp_126 & (mux_218_nl) & and_208_cse & and_dcpl_160 &
      (else_7_else_1_else_div_5cyc_st_3[0]);
  assign mux_219_cse = MUX_s_1_2_2({(~(or_cse | (~ and_tmp_107))) , and_tmp_107},
      or_tmp_652);
  assign mux_226_nl = MUX_s_1_2_2({(~(or_cse | (~ mux_tmp_170))) , mux_tmp_170},
      or_tmp_689);
  assign and_1449_cse = or_tmp_126 & (mux_226_nl) & and_208_cse & (~ (else_7_else_1_else_div_5cyc_st_3[1]))
      & (else_7_else_1_else_div_5cyc_st_3[2]) & (~ (else_7_else_1_else_div_5cyc_st_3[0]));
  assign mux_229_cse = MUX_s_1_2_2({(~(or_cse | (~ mux_228_cse))) , mux_228_cse},
      or_tmp_689);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      V_OUT_rsc_mgc_out_stdreg_d <= 10'b0;
      S_OUT_rsc_mgc_out_stdreg_d <= 10'b0;
      H_OUT_rsc_mgc_out_stdreg_d <= 10'b0;
      else_7_acc_1_psp_sg1_sva <= 11'b0;
      h_4_sva_duc <= 18'b0;
      else_7_if_1_div_5cyc_st_5 <= 3'b0;
      h_6_sva_duc <= 18'b0;
      h_5_sva_duc <= 18'b0;
      else_7_else_1_if_div_5cyc_st_5 <= 3'b0;
      else_7_else_1_else_div_5cyc_st_5 <= 3'b0;
      else_7_else_1_equal_svs_st_5 <= 1'b0;
      else_7_and_5_itm_5 <= 1'b0;
      else_7_equal_svs_5 <= 1'b0;
      else_7_else_1_equal_svs_5 <= 1'b0;
      else_7_equal_svs_st_5 <= 1'b0;
      acc_5_itm_5 <= 9'b0;
      acc_4_itm_2 <= 10'b0;
      unequal_tmp_6 <= 1'b0;
      acc_2_psp_sva_st_5 <= 10'b0;
      mut_62_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_12_sg1 <= 10'b0;
      mut_66_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_16_sg1 <= 10'b0;
      mut_70_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_20_sg1 <= 10'b0;
      mut_74_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_24_sg1 <= 10'b0;
      mut_18_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_8_sg1 <= 10'b0;
      else_7_if_1_div_5cyc_st_4 <= 3'b0;
      mut_42_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_8_sg1 <= 10'b0;
      mut_46_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_12_sg1 <= 10'b0;
      mut_50_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_16_sg1 <= 10'b0;
      mut_54_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_20_sg1 <= 10'b0;
      mut_58_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_24_sg1 <= 10'b0;
      else_7_else_1_if_div_5cyc_st_4 <= 3'b0;
      mut_22_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_8_sg1 <= 10'b0;
      mut_26_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_12_sg1 <= 10'b0;
      mut_30_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_16_sg1 <= 10'b0;
      mut_34_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_20_sg1 <= 10'b0;
      mut_38_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_24_sg1 <= 10'b0;
      else_7_else_1_else_div_5cyc_st_4 <= 3'b0;
      else_7_else_1_equal_svs_st_4 <= 1'b0;
      else_7_equal_svs_st_4 <= 1'b0;
      acc_2_psp_sva_st_4 <= 10'b0;
      else_7_if_div_2cyc_st_3 <= 1'b0;
      mut_61_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_11_sg1 <= 10'b0;
      mut_65_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_15_sg1 <= 10'b0;
      mut_69_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_19_sg1 <= 10'b0;
      mut_73_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_23_sg1 <= 10'b0;
      mut_17_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_7_sg1 <= 10'b0;
      else_7_if_1_div_5cyc_st_3 <= 3'b0;
      mut_41_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_7_sg1 <= 10'b0;
      mut_45_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_11_sg1 <= 10'b0;
      mut_49_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_15_sg1 <= 10'b0;
      mut_53_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_19_sg1 <= 10'b0;
      mut_57_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_23_sg1 <= 10'b0;
      else_7_else_1_if_div_5cyc_st_3 <= 3'b0;
      mut_21_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_7_sg1 <= 10'b0;
      mut_25_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_11_sg1 <= 10'b0;
      mut_29_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_15_sg1 <= 10'b0;
      mut_33_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_19_sg1 <= 10'b0;
      mut_37_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_23_sg1 <= 10'b0;
      else_7_else_1_else_div_5cyc_st_3 <= 3'b0;
      else_7_else_1_equal_svs_st_3 <= 1'b0;
      else_7_equal_svs_st_3 <= 1'b0;
      max_sg1_lpi_dfm_3_st_3 <= 10'b0;
      acc_2_psp_sva_st_3 <= 10'b0;
      mut_60_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_10_sg1 <= 10'b0;
      mut_64_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_14_sg1 <= 10'b0;
      mut_68_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_18_sg1 <= 10'b0;
      mut_72_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_22_sg1 <= 10'b0;
      mut_16_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_6_sg1 <= 10'b0;
      else_7_if_1_div_5cyc_st_2 <= 3'b0;
      mut_40_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_6_sg1 <= 10'b0;
      mut_44_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_10_sg1 <= 10'b0;
      mut_48_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_14_sg1 <= 10'b0;
      mut_52_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_18_sg1 <= 10'b0;
      mut_56_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_22_sg1 <= 10'b0;
      else_7_else_1_if_div_5cyc_st_2 <= 3'b0;
      mut_20_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_6_sg1 <= 10'b0;
      mut_24_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_10_sg1 <= 10'b0;
      mut_28_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_14_sg1 <= 10'b0;
      mut_32_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_18_sg1 <= 10'b0;
      mut_36_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_22_sg1 <= 10'b0;
      else_7_else_1_else_div_5cyc_st_2 <= 3'b0;
      else_7_else_1_equal_svs_st_2 <= 1'b0;
      else_7_equal_svs_st_2 <= 1'b0;
      acc_2_psp_sva_st_2 <= 10'b0;
      reg_div_mgc_div_16_b_cse <= 10'b0;
      reg_div_mgc_div_15_b_cse <= 10'b0;
      else_7_if_div_2cyc_st_1 <= 1'b0;
      mut_59_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_9_sg1 <= 10'b0;
      mut_63_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_13_sg1 <= 10'b0;
      mut_67_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_17_sg1 <= 10'b0;
      mut_71_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_21_sg1 <= 10'b0;
      mut_15_sg1 <= 10'b0;
      else_7_if_1_conc_1_tmp_mut_5_sg1 <= 10'b0;
      else_7_if_1_div_5cyc_st_1 <= 3'b0;
      mut_39_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_5_sg1 <= 10'b0;
      mut_43_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_9_sg1 <= 10'b0;
      mut_47_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_13_sg1 <= 10'b0;
      mut_51_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_17_sg1 <= 10'b0;
      mut_55_sg1 <= 10'b0;
      else_7_else_1_if_conc_1_tmp_mut_21_sg1 <= 10'b0;
      else_7_else_1_if_div_5cyc_st_1 <= 3'b0;
      mut_19_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_5_sg1 <= 10'b0;
      mut_23_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_9_sg1 <= 10'b0;
      mut_27_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_13_sg1 <= 10'b0;
      mut_31_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_17_sg1 <= 10'b0;
      mut_35_sg1 <= 10'b0;
      else_7_else_1_else_conc_1_tmp_mut_21_sg1 <= 10'b0;
      else_7_else_1_else_div_5cyc_st_1 <= 3'b0;
      else_7_else_1_equal_svs_st_1 <= 1'b0;
      else_7_equal_svs_st_1 <= 1'b0;
      reg_max_sg1_lpi_dfm_3_st_1_cse <= 10'b0;
      acc_2_psp_sva_st_1 <= 10'b0;
      else_7_if_div_2cyc <= 1'b0;
      else_7_if_1_div_5cyc <= 3'b0;
      else_7_else_1_if_div_5cyc <= 3'b0;
      else_7_else_1_else_div_5cyc <= 3'b0;
      else_7_equal_svs <= 1'b0;
      unequal_tmp_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      else_7_if_conc_1_tmp_mut_1_sg1 <= 10'b0;
      else_7_if_conc_1_tmp_mut_sg1 <= 10'b0;
      else_7_if_div_2cyc_st_2 <= 1'b0;
      max_sg1_lpi_dfm_3_st_2 <= 10'b0;
      acc_5_itm_4 <= 9'b0;
      acc_4_itm_1 <= 10'b0;
      else_7_and_5_itm_4 <= 1'b0;
      else_7_equal_svs_4 <= 1'b0;
      unequal_tmp_5 <= 1'b0;
      else_7_else_1_equal_svs_4 <= 1'b0;
      s_sg1_1_sva_2_duc <= 18'b0;
      unequal_tmp_9 <= 1'b0;
      unequal_tmp_4 <= 1'b0;
      acc_5_itm_3 <= 9'b0;
      else_7_and_5_itm_3 <= 1'b0;
      else_7_equal_svs_3 <= 1'b0;
      else_7_else_1_equal_svs_3 <= 1'b0;
      acc_5_itm_2 <= 9'b0;
      else_7_and_5_itm_2 <= 1'b0;
      else_7_equal_svs_2 <= 1'b0;
      unequal_tmp_8 <= 1'b0;
      unequal_tmp_3 <= 1'b0;
      else_7_else_1_equal_svs_2 <= 1'b0;
      acc_5_itm_1 <= 9'b0;
      else_7_and_5_itm_1 <= 1'b0;
      unequal_tmp_2 <= 1'b0;
      else_7_else_1_equal_svs_1 <= 1'b0;
      reg_div_mgc_div_11_b_tmp <= 10'b0;
      reg_div_mgc_div_11_a_tmp <= 10'b0;
      reg_div_mgc_div_12_b_tmp <= 10'b0;
      reg_div_mgc_div_12_a_tmp <= 10'b0;
      reg_div_mgc_div_13_b_tmp <= 10'b0;
      reg_div_mgc_div_13_a_tmp <= 10'b0;
      reg_div_mgc_div_14_b_tmp <= 10'b0;
      reg_div_mgc_div_14_a_tmp <= 10'b0;
      reg_div_mgc_div_b_tmp <= 10'b0;
      reg_div_mgc_div_a_tmp <= 10'b0;
      reg_div_mgc_div_6_b_tmp <= 10'b0;
      reg_div_mgc_div_6_a_tmp <= 10'b0;
      reg_div_mgc_div_7_b_tmp <= 10'b0;
      reg_div_mgc_div_7_a_tmp <= 10'b0;
      reg_div_mgc_div_8_b_tmp <= 10'b0;
      reg_div_mgc_div_8_a_tmp <= 10'b0;
      reg_div_mgc_div_9_b_tmp <= 10'b0;
      reg_div_mgc_div_9_a_tmp <= 10'b0;
      reg_div_mgc_div_10_b_tmp <= 10'b0;
      reg_div_mgc_div_10_a_tmp <= 10'b0;
      reg_div_mgc_div_1_b_tmp <= 10'b0;
      reg_div_mgc_div_1_a_tmp <= 10'b0;
      reg_div_mgc_div_2_b_tmp <= 10'b0;
      reg_div_mgc_div_2_a_tmp <= 10'b0;
      reg_div_mgc_div_3_b_tmp <= 10'b0;
      reg_div_mgc_div_3_a_tmp <= 10'b0;
      reg_div_mgc_div_4_b_tmp <= 10'b0;
      reg_div_mgc_div_4_a_tmp <= 10'b0;
      reg_div_mgc_div_5_b_tmp <= 10'b0;
      reg_div_mgc_div_5_a_tmp <= 10'b0;
    end
    else begin
      V_OUT_rsc_mgc_out_stdreg_d <= MUX_v_10_2_2({V_OUT_rsc_mgc_out_stdreg_d , ({1'b0
          , acc_5_itm_5})}, main_stage_0_6);
      S_OUT_rsc_mgc_out_stdreg_d <= MUX_v_10_2_2({S_OUT_rsc_mgc_out_stdreg_d , acc_4_itm_2},
          main_stage_0_6);
      H_OUT_rsc_mgc_out_stdreg_d <= MUX_v_10_2_2({H_OUT_rsc_mgc_out_stdreg_d , (({((MUX_v_7_2_2({(else_7_acc_1_psp_sg1_sva_1[10:4])
          , (({1'b1 , (else_7_acc_1_itm[16:11])}) + 7'b101101)}, else_7_acc_1_psp_sg1_sva_1[10]))
          & ({{6{unequal_tmp_6}}, unequal_tmp_6})) , (h_1_sg1_lpi_dfm_1[3:1])}) +
          conv_u2u_1_10(h_1_sg1_lpi_dfm_1[0]))}, main_stage_0_6);
      else_7_acc_1_psp_sg1_sva <= MUX_v_11_2_2({else_7_acc_1_psp_sg1_sva , (else_7_acc_1_itm[17:7])},
          (~ and_1892_cse) & main_stage_0_6);
      h_4_sva_duc <= MUX1HOT_v_18_6_2({(div_mgc_div_11_z[17:0]) , (div_mgc_div_12_z[17:0])
          , (div_mgc_div_13_z[17:0]) , (div_mgc_div_14_z[17:0]) , (div_mgc_div_z[17:0])
          , h_4_sva_duc}, {(or_489_cse & and_dcpl_521 & and_dcpl_503) , (or_489_cse
          & and_dcpl_521 & and_dcpl_506) , (or_489_cse & and_dcpl_531 & and_dcpl_503)
          , (or_489_cse & and_dcpl_531 & and_dcpl_506) , (or_489_cse & and_dcpl_521
          & and_dcpl_515) , (and_1892_cse | and_dcpl_518 | (~(main_stage_0_6 & else_7_equal_svs_st_5)))});
      else_7_if_1_div_5cyc_st_5 <= else_7_if_1_div_5cyc_st_4;
      h_6_sva_duc <= MUX1HOT_v_18_6_2({(div_mgc_div_6_z[17:0]) , (div_mgc_div_7_z[17:0])
          , (div_mgc_div_8_z[17:0]) , (div_mgc_div_9_z[17:0]) , (div_mgc_div_10_z[17:0])
          , h_6_sva_duc}, {(or_489_cse & and_dcpl_589 & and_588_cse) , (or_489_cse
          & and_dcpl_589 & and_590_cse) , (or_489_cse & and_dcpl_589 & and_592_cse)
          , (or_489_cse & and_dcpl_589 & and_594_cse) , (or_489_cse & and_dcpl_589
          & and_596_cse) , (and_1892_cse | or_dcpl_462 | (~ else_7_else_1_equal_svs_st_5)
          | and_dcpl_574)});
      h_5_sva_duc <= MUX1HOT_v_18_6_2({(div_mgc_div_1_z[17:0]) , (div_mgc_div_2_z[17:0])
          , (div_mgc_div_3_z[17:0]) , (div_mgc_div_4_z[17:0]) , (div_mgc_div_5_z[17:0])
          , h_5_sva_duc}, {(or_489_cse & and_dcpl_661 & and_660_cse) , (or_489_cse
          & and_dcpl_661 & and_662_cse) , (or_489_cse & and_dcpl_661 & and_664_cse)
          , (or_489_cse & and_dcpl_661 & and_666_cse) , (or_489_cse & and_dcpl_661
          & and_668_cse) , (and_1892_cse | or_dcpl_462 | else_7_else_1_equal_svs_st_5
          | and_dcpl_646)});
      else_7_else_1_if_div_5cyc_st_5 <= else_7_else_1_if_div_5cyc_st_4;
      else_7_else_1_else_div_5cyc_st_5 <= else_7_else_1_else_div_5cyc_st_4;
      else_7_else_1_equal_svs_st_5 <= else_7_else_1_equal_svs_st_4;
      else_7_and_5_itm_5 <= else_7_and_5_itm_4;
      else_7_equal_svs_5 <= else_7_equal_svs_4;
      else_7_else_1_equal_svs_5 <= else_7_else_1_equal_svs_4;
      else_7_equal_svs_st_5 <= else_7_equal_svs_st_4;
      acc_5_itm_5 <= acc_5_itm_4;
      acc_4_itm_2 <= acc_4_itm_1;
      unequal_tmp_6 <= unequal_tmp_5;
      acc_2_psp_sva_st_5 <= acc_2_psp_sva_st_4;
      mut_62_sg1 <= mut_61_sg1;
      else_7_if_1_conc_1_tmp_mut_12_sg1 <= else_7_if_1_conc_1_tmp_mut_11_sg1;
      mut_66_sg1 <= mut_65_sg1;
      else_7_if_1_conc_1_tmp_mut_16_sg1 <= else_7_if_1_conc_1_tmp_mut_15_sg1;
      mut_70_sg1 <= mut_69_sg1;
      else_7_if_1_conc_1_tmp_mut_20_sg1 <= else_7_if_1_conc_1_tmp_mut_19_sg1;
      mut_74_sg1 <= mut_73_sg1;
      else_7_if_1_conc_1_tmp_mut_24_sg1 <= else_7_if_1_conc_1_tmp_mut_23_sg1;
      mut_18_sg1 <= mut_17_sg1;
      else_7_if_1_conc_1_tmp_mut_8_sg1 <= else_7_if_1_conc_1_tmp_mut_7_sg1;
      else_7_if_1_div_5cyc_st_4 <= else_7_if_1_div_5cyc_st_3;
      mut_42_sg1 <= mut_41_sg1;
      else_7_else_1_if_conc_1_tmp_mut_8_sg1 <= else_7_else_1_if_conc_1_tmp_mut_7_sg1;
      mut_46_sg1 <= mut_45_sg1;
      else_7_else_1_if_conc_1_tmp_mut_12_sg1 <= else_7_else_1_if_conc_1_tmp_mut_11_sg1;
      mut_50_sg1 <= mut_49_sg1;
      else_7_else_1_if_conc_1_tmp_mut_16_sg1 <= else_7_else_1_if_conc_1_tmp_mut_15_sg1;
      mut_54_sg1 <= mut_53_sg1;
      else_7_else_1_if_conc_1_tmp_mut_20_sg1 <= else_7_else_1_if_conc_1_tmp_mut_19_sg1;
      mut_58_sg1 <= mut_57_sg1;
      else_7_else_1_if_conc_1_tmp_mut_24_sg1 <= else_7_else_1_if_conc_1_tmp_mut_23_sg1;
      else_7_else_1_if_div_5cyc_st_4 <= else_7_else_1_if_div_5cyc_st_3;
      mut_22_sg1 <= mut_21_sg1;
      else_7_else_1_else_conc_1_tmp_mut_8_sg1 <= else_7_else_1_else_conc_1_tmp_mut_7_sg1;
      mut_26_sg1 <= mut_25_sg1;
      else_7_else_1_else_conc_1_tmp_mut_12_sg1 <= else_7_else_1_else_conc_1_tmp_mut_11_sg1;
      mut_30_sg1 <= mut_29_sg1;
      else_7_else_1_else_conc_1_tmp_mut_16_sg1 <= else_7_else_1_else_conc_1_tmp_mut_15_sg1;
      mut_34_sg1 <= mut_33_sg1;
      else_7_else_1_else_conc_1_tmp_mut_20_sg1 <= else_7_else_1_else_conc_1_tmp_mut_19_sg1;
      mut_38_sg1 <= mut_37_sg1;
      else_7_else_1_else_conc_1_tmp_mut_24_sg1 <= else_7_else_1_else_conc_1_tmp_mut_23_sg1;
      else_7_else_1_else_div_5cyc_st_4 <= else_7_else_1_else_div_5cyc_st_3;
      else_7_else_1_equal_svs_st_4 <= else_7_else_1_equal_svs_st_3;
      else_7_equal_svs_st_4 <= else_7_equal_svs_st_3;
      acc_2_psp_sva_st_4 <= acc_2_psp_sva_st_3;
      else_7_if_div_2cyc_st_3 <= else_7_if_div_2cyc_st_2;
      mut_61_sg1 <= mut_60_sg1;
      else_7_if_1_conc_1_tmp_mut_11_sg1 <= else_7_if_1_conc_1_tmp_mut_10_sg1;
      mut_65_sg1 <= mut_64_sg1;
      else_7_if_1_conc_1_tmp_mut_15_sg1 <= else_7_if_1_conc_1_tmp_mut_14_sg1;
      mut_69_sg1 <= mut_68_sg1;
      else_7_if_1_conc_1_tmp_mut_19_sg1 <= else_7_if_1_conc_1_tmp_mut_18_sg1;
      mut_73_sg1 <= mut_72_sg1;
      else_7_if_1_conc_1_tmp_mut_23_sg1 <= else_7_if_1_conc_1_tmp_mut_22_sg1;
      mut_17_sg1 <= mut_16_sg1;
      else_7_if_1_conc_1_tmp_mut_7_sg1 <= else_7_if_1_conc_1_tmp_mut_6_sg1;
      else_7_if_1_div_5cyc_st_3 <= else_7_if_1_div_5cyc_st_2;
      mut_41_sg1 <= mut_40_sg1;
      else_7_else_1_if_conc_1_tmp_mut_7_sg1 <= else_7_else_1_if_conc_1_tmp_mut_6_sg1;
      mut_45_sg1 <= mut_44_sg1;
      else_7_else_1_if_conc_1_tmp_mut_11_sg1 <= else_7_else_1_if_conc_1_tmp_mut_10_sg1;
      mut_49_sg1 <= mut_48_sg1;
      else_7_else_1_if_conc_1_tmp_mut_15_sg1 <= else_7_else_1_if_conc_1_tmp_mut_14_sg1;
      mut_53_sg1 <= mut_52_sg1;
      else_7_else_1_if_conc_1_tmp_mut_19_sg1 <= else_7_else_1_if_conc_1_tmp_mut_18_sg1;
      mut_57_sg1 <= mut_56_sg1;
      else_7_else_1_if_conc_1_tmp_mut_23_sg1 <= else_7_else_1_if_conc_1_tmp_mut_22_sg1;
      else_7_else_1_if_div_5cyc_st_3 <= else_7_else_1_if_div_5cyc_st_2;
      mut_21_sg1 <= mut_20_sg1;
      else_7_else_1_else_conc_1_tmp_mut_7_sg1 <= else_7_else_1_else_conc_1_tmp_mut_6_sg1;
      mut_25_sg1 <= mut_24_sg1;
      else_7_else_1_else_conc_1_tmp_mut_11_sg1 <= else_7_else_1_else_conc_1_tmp_mut_10_sg1;
      mut_29_sg1 <= mut_28_sg1;
      else_7_else_1_else_conc_1_tmp_mut_15_sg1 <= else_7_else_1_else_conc_1_tmp_mut_14_sg1;
      mut_33_sg1 <= mut_32_sg1;
      else_7_else_1_else_conc_1_tmp_mut_19_sg1 <= else_7_else_1_else_conc_1_tmp_mut_18_sg1;
      mut_37_sg1 <= mut_36_sg1;
      else_7_else_1_else_conc_1_tmp_mut_23_sg1 <= else_7_else_1_else_conc_1_tmp_mut_22_sg1;
      else_7_else_1_else_div_5cyc_st_3 <= else_7_else_1_else_div_5cyc_st_2;
      else_7_else_1_equal_svs_st_3 <= else_7_else_1_equal_svs_st_2;
      else_7_equal_svs_st_3 <= else_7_equal_svs_st_2;
      max_sg1_lpi_dfm_3_st_3 <= max_sg1_lpi_dfm_3_st_2;
      acc_2_psp_sva_st_3 <= acc_2_psp_sva_st_2;
      mut_60_sg1 <= mut_59_sg1;
      else_7_if_1_conc_1_tmp_mut_10_sg1 <= else_7_if_1_conc_1_tmp_mut_9_sg1;
      mut_64_sg1 <= mut_63_sg1;
      else_7_if_1_conc_1_tmp_mut_14_sg1 <= else_7_if_1_conc_1_tmp_mut_13_sg1;
      mut_68_sg1 <= mut_67_sg1;
      else_7_if_1_conc_1_tmp_mut_18_sg1 <= else_7_if_1_conc_1_tmp_mut_17_sg1;
      mut_72_sg1 <= mut_71_sg1;
      else_7_if_1_conc_1_tmp_mut_22_sg1 <= else_7_if_1_conc_1_tmp_mut_21_sg1;
      mut_16_sg1 <= mut_15_sg1;
      else_7_if_1_conc_1_tmp_mut_6_sg1 <= else_7_if_1_conc_1_tmp_mut_5_sg1;
      else_7_if_1_div_5cyc_st_2 <= else_7_if_1_div_5cyc_st_1;
      mut_40_sg1 <= mut_39_sg1;
      else_7_else_1_if_conc_1_tmp_mut_6_sg1 <= else_7_else_1_if_conc_1_tmp_mut_5_sg1;
      mut_44_sg1 <= mut_43_sg1;
      else_7_else_1_if_conc_1_tmp_mut_10_sg1 <= else_7_else_1_if_conc_1_tmp_mut_9_sg1;
      mut_48_sg1 <= mut_47_sg1;
      else_7_else_1_if_conc_1_tmp_mut_14_sg1 <= else_7_else_1_if_conc_1_tmp_mut_13_sg1;
      mut_52_sg1 <= mut_51_sg1;
      else_7_else_1_if_conc_1_tmp_mut_18_sg1 <= else_7_else_1_if_conc_1_tmp_mut_17_sg1;
      mut_56_sg1 <= mut_55_sg1;
      else_7_else_1_if_conc_1_tmp_mut_22_sg1 <= else_7_else_1_if_conc_1_tmp_mut_21_sg1;
      else_7_else_1_if_div_5cyc_st_2 <= else_7_else_1_if_div_5cyc_st_1;
      mut_20_sg1 <= mut_19_sg1;
      else_7_else_1_else_conc_1_tmp_mut_6_sg1 <= else_7_else_1_else_conc_1_tmp_mut_5_sg1;
      mut_24_sg1 <= mut_23_sg1;
      else_7_else_1_else_conc_1_tmp_mut_10_sg1 <= else_7_else_1_else_conc_1_tmp_mut_9_sg1;
      mut_28_sg1 <= mut_27_sg1;
      else_7_else_1_else_conc_1_tmp_mut_14_sg1 <= else_7_else_1_else_conc_1_tmp_mut_13_sg1;
      mut_32_sg1 <= mut_31_sg1;
      else_7_else_1_else_conc_1_tmp_mut_18_sg1 <= else_7_else_1_else_conc_1_tmp_mut_17_sg1;
      mut_36_sg1 <= mut_35_sg1;
      else_7_else_1_else_conc_1_tmp_mut_22_sg1 <= else_7_else_1_else_conc_1_tmp_mut_21_sg1;
      else_7_else_1_else_div_5cyc_st_2 <= else_7_else_1_else_div_5cyc_st_1;
      else_7_else_1_equal_svs_st_2 <= else_7_else_1_equal_svs_st_1;
      else_7_equal_svs_st_2 <= else_7_equal_svs_st_1;
      acc_2_psp_sva_st_2 <= acc_2_psp_sva_st_1;
      reg_div_mgc_div_16_b_cse <= MUX_v_10_2_2({mux1h_38_tmp , reg_div_mgc_div_16_b_cse},
          or_dcpl_790);
      reg_div_mgc_div_15_b_cse <= MUX_v_10_2_2({mux1h_38_tmp , reg_div_mgc_div_15_b_cse},
          or_dcpl_792);
      else_7_if_div_2cyc_st_1 <= MUX_s_1_2_2({(~ else_7_if_div_2cyc) , else_7_if_div_2cyc_st_1},
          not_tmp_349);
      mut_59_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_59_sg1}, and_1483_cse);
      else_7_if_1_conc_1_tmp_mut_9_sg1 <= MUX_v_10_2_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_9_sg1}, and_1483_cse);
      mut_63_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_63_sg1}, and_1483_cse);
      else_7_if_1_conc_1_tmp_mut_13_sg1 <= MUX_v_10_2_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_13_sg1}, and_1483_cse);
      mut_67_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_67_sg1}, and_1483_cse);
      else_7_if_1_conc_1_tmp_mut_17_sg1 <= MUX_v_10_2_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_17_sg1}, and_1483_cse);
      mut_71_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_71_sg1}, and_1483_cse);
      else_7_if_1_conc_1_tmp_mut_21_sg1 <= MUX_v_10_2_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_21_sg1}, and_1483_cse);
      mut_15_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_15_sg1}, and_1483_cse);
      else_7_if_1_conc_1_tmp_mut_5_sg1 <= MUX_v_10_2_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_5_sg1}, and_1483_cse);
      else_7_if_1_div_5cyc_st_1 <= MUX_v_3_2_2({else_7_if_1_acc_tmp , else_7_if_1_div_5cyc_st_1},
          and_1483_cse);
      mut_39_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_39_sg1}, and_1483_cse);
      else_7_else_1_if_conc_1_tmp_mut_5_sg1 <= MUX_v_10_2_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_5_sg1}, and_1483_cse);
      mut_43_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_43_sg1}, and_1483_cse);
      else_7_else_1_if_conc_1_tmp_mut_9_sg1 <= MUX_v_10_2_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_9_sg1}, and_1483_cse);
      mut_47_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_47_sg1}, and_1483_cse);
      else_7_else_1_if_conc_1_tmp_mut_13_sg1 <= MUX_v_10_2_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_13_sg1}, and_1483_cse);
      mut_51_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_51_sg1}, and_1483_cse);
      else_7_else_1_if_conc_1_tmp_mut_17_sg1 <= MUX_v_10_2_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_17_sg1}, and_1483_cse);
      mut_55_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_55_sg1}, and_1483_cse);
      else_7_else_1_if_conc_1_tmp_mut_21_sg1 <= MUX_v_10_2_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_21_sg1}, and_1483_cse);
      else_7_else_1_if_div_5cyc_st_1 <= MUX_v_3_2_2({else_7_else_1_if_acc_tmp , else_7_else_1_if_div_5cyc_st_1},
          and_1483_cse);
      mut_19_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_19_sg1}, and_1483_cse);
      else_7_else_1_else_conc_1_tmp_mut_5_sg1 <= MUX_v_10_2_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_5_sg1}, and_1483_cse);
      mut_23_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_23_sg1}, and_1483_cse);
      else_7_else_1_else_conc_1_tmp_mut_9_sg1 <= MUX_v_10_2_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_9_sg1}, and_1483_cse);
      mut_27_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_27_sg1}, and_1483_cse);
      else_7_else_1_else_conc_1_tmp_mut_13_sg1 <= MUX_v_10_2_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_13_sg1}, and_1483_cse);
      mut_31_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_31_sg1}, and_1483_cse);
      else_7_else_1_else_conc_1_tmp_mut_17_sg1 <= MUX_v_10_2_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_17_sg1}, and_1483_cse);
      mut_35_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , mut_35_sg1}, and_1483_cse);
      else_7_else_1_else_conc_1_tmp_mut_21_sg1 <= MUX_v_10_2_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_21_sg1}, and_1483_cse);
      else_7_else_1_else_div_5cyc_st_1 <= MUX_v_3_2_2({else_7_else_1_else_acc_tmp
          , else_7_else_1_else_div_5cyc_st_1}, and_1483_cse);
      else_7_else_1_equal_svs_st_1 <= MUX_s_1_2_2({else_7_else_1_equal_tmp , else_7_else_1_equal_svs_st_1},
          and_1483_cse);
      else_7_equal_svs_st_1 <= MUX_s_1_2_2({else_7_equal_tmp , else_7_equal_svs_st_1},
          and_1483_cse);
      reg_max_sg1_lpi_dfm_3_st_1_cse <= MUX_v_10_2_2({mux1h_38_tmp , reg_max_sg1_lpi_dfm_3_st_1_cse},
          and_1483_cse);
      acc_2_psp_sva_st_1 <= acc_itm[10:1];
      else_7_if_div_2cyc <= MUX_s_1_2_2({(~ else_7_if_div_2cyc) , else_7_if_div_2cyc},
          not_tmp_349);
      else_7_if_1_div_5cyc <= MUX_v_3_2_2({else_7_if_1_acc_tmp , else_7_if_1_div_5cyc},
          ~((~(and_dcpl_1354 & and_dcpl_1352 & and_dcpl_1350 & and_dcpl_1348)) &
          else_7_equal_tmp));
      else_7_else_1_if_div_5cyc <= MUX_v_3_2_2({else_7_else_1_if_acc_tmp , else_7_else_1_if_div_5cyc},
          and_1483_cse | else_7_equal_tmp | (~ else_7_else_1_equal_tmp));
      else_7_else_1_else_div_5cyc <= MUX_v_3_2_2({else_7_else_1_else_acc_tmp , else_7_else_1_else_div_5cyc},
          and_1483_cse | else_7_equal_tmp | else_7_else_1_equal_tmp);
      else_7_equal_svs <= MUX_s_1_2_2({else_7_equal_tmp , else_7_equal_svs}, and_1483_cse);
      unequal_tmp_1 <= MUX_s_1_2_2({unequal_tmp_10 , unequal_tmp_1}, and_1483_cse);
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      else_7_if_conc_1_tmp_mut_1_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , else_7_if_conc_1_tmp_mut_1_sg1},
          or_dcpl_790);
      else_7_if_conc_1_tmp_mut_sg1 <= MUX_v_10_2_2({(acc_itm[10:1]) , else_7_if_conc_1_tmp_mut_sg1},
          or_dcpl_792);
      else_7_if_div_2cyc_st_2 <= else_7_if_div_2cyc_st_1;
      max_sg1_lpi_dfm_3_st_2 <= reg_max_sg1_lpi_dfm_3_st_1_cse;
      acc_5_itm_4 <= acc_5_itm_3;
      acc_4_itm_1 <= nl_acc_4_itm_1[9:0];
      else_7_and_5_itm_4 <= else_7_and_5_itm_3;
      else_7_equal_svs_4 <= else_7_equal_svs_3;
      unequal_tmp_5 <= unequal_tmp_4;
      else_7_else_1_equal_svs_4 <= else_7_else_1_equal_svs_3;
      s_sg1_1_sva_2_duc <= MUX1HOT_v_18_3_2({(div_mgc_div_16_z_oreg[17:0]) , (div_mgc_div_15_z_oreg[17:0])
          , s_sg1_1_sva_2_duc}, {(and_tmp_116 & main_stage_0_4 & (~ else_7_if_div_2cyc_st_3))
          , (and_tmp_116 & main_stage_0_4 & else_7_if_div_2cyc_st_3) , (~(and_tmp_116
          & main_stage_0_4))});
      unequal_tmp_9 <= unequal_tmp_8;
      unequal_tmp_4 <= unequal_tmp_3;
      acc_5_itm_3 <= acc_5_itm_2;
      else_7_and_5_itm_3 <= else_7_and_5_itm_2;
      else_7_equal_svs_3 <= else_7_equal_svs_2;
      else_7_else_1_equal_svs_3 <= else_7_else_1_equal_svs_2;
      acc_5_itm_2 <= acc_5_itm_1;
      else_7_and_5_itm_2 <= else_7_and_5_itm_1;
      else_7_equal_svs_2 <= else_7_equal_svs;
      unequal_tmp_8 <= unequal_tmp_1;
      unequal_tmp_3 <= unequal_tmp_2;
      else_7_else_1_equal_svs_2 <= else_7_else_1_equal_svs_1;
      acc_5_itm_1 <= nl_acc_5_itm_1[8:0];
      else_7_and_5_itm_1 <= MUX_s_1_2_2({(else_7_else_1_equal_tmp & (~ else_7_equal_tmp))
          , else_7_and_5_itm_1}, and_1483_cse);
      unequal_tmp_2 <= or_cse;
      else_7_else_1_equal_svs_1 <= else_7_else_1_equal_tmp;
      reg_div_mgc_div_11_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_59_sg1
          , mut_60_sg1 , mut_61_sg1 , mut_62_sg1}, {and_713_cse , and_718_cse , and_723_cse
          , and_730_cse , mux_95_cse});
      reg_div_mgc_div_11_a_tmp <= MUX1HOT_v_10_5_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_9_sg1 , else_7_if_1_conc_1_tmp_mut_10_sg1
          , else_7_if_1_conc_1_tmp_mut_11_sg1 , else_7_if_1_conc_1_tmp_mut_12_sg1},
          {and_713_cse , and_718_cse , and_723_cse , and_730_cse , mux_95_cse});
      reg_div_mgc_div_12_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_63_sg1
          , mut_64_sg1 , mut_65_sg1 , mut_66_sg1}, {and_759_cse , and_764_cse , and_769_cse
          , and_776_cse , mux_106_cse});
      reg_div_mgc_div_12_a_tmp <= MUX1HOT_v_10_5_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_13_sg1 , else_7_if_1_conc_1_tmp_mut_14_sg1
          , else_7_if_1_conc_1_tmp_mut_15_sg1 , else_7_if_1_conc_1_tmp_mut_16_sg1},
          {and_759_cse , and_764_cse , and_769_cse , and_776_cse , mux_106_cse});
      reg_div_mgc_div_13_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_67_sg1
          , mut_68_sg1 , mut_69_sg1 , mut_70_sg1}, {and_805_cse , and_810_cse , and_815_cse
          , and_822_cse , mux_117_cse});
      reg_div_mgc_div_13_a_tmp <= MUX1HOT_v_10_5_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_17_sg1 , else_7_if_1_conc_1_tmp_mut_18_sg1
          , else_7_if_1_conc_1_tmp_mut_19_sg1 , else_7_if_1_conc_1_tmp_mut_20_sg1},
          {and_805_cse , and_810_cse , and_815_cse , and_822_cse , mux_117_cse});
      reg_div_mgc_div_14_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_71_sg1
          , mut_72_sg1 , mut_73_sg1 , mut_74_sg1}, {and_851_cse , and_856_cse , and_861_cse
          , and_868_cse , mux_128_cse});
      reg_div_mgc_div_14_a_tmp <= MUX1HOT_v_10_5_2({(else_7_if_1_acc_1_itm[10:1])
          , else_7_if_1_conc_1_tmp_mut_21_sg1 , else_7_if_1_conc_1_tmp_mut_22_sg1
          , else_7_if_1_conc_1_tmp_mut_23_sg1 , else_7_if_1_conc_1_tmp_mut_24_sg1},
          {and_851_cse , and_856_cse , and_861_cse , and_868_cse , mux_128_cse});
      reg_div_mgc_div_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_15_sg1 , mut_16_sg1
          , mut_17_sg1 , mut_18_sg1}, {and_897_cse , and_902_cse , and_907_cse ,
          and_913_cse , mux_145_cse});
      reg_div_mgc_div_a_tmp <= MUX1HOT_v_10_5_2({(else_7_if_1_acc_1_itm[10:1]) ,
          else_7_if_1_conc_1_tmp_mut_5_sg1 , else_7_if_1_conc_1_tmp_mut_6_sg1 , else_7_if_1_conc_1_tmp_mut_7_sg1
          , else_7_if_1_conc_1_tmp_mut_8_sg1}, {and_897_cse , and_902_cse , and_907_cse
          , and_913_cse , mux_145_cse});
      reg_div_mgc_div_6_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_39_sg1 ,
          mut_40_sg1 , mut_41_sg1 , mut_42_sg1}, {and_938_cse , and_945_cse , and_952_cse
          , and_960_cse , mux_157_cse});
      reg_div_mgc_div_6_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_5_sg1 , else_7_else_1_if_conc_1_tmp_mut_6_sg1
          , else_7_else_1_if_conc_1_tmp_mut_7_sg1 , else_7_else_1_if_conc_1_tmp_mut_8_sg1},
          {and_938_cse , and_945_cse , and_952_cse , and_960_cse , mux_157_cse});
      reg_div_mgc_div_7_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_43_sg1 ,
          mut_44_sg1 , mut_45_sg1 , mut_46_sg1}, {and_994_cse , and_1000_cse , and_1007_cse
          , and_1015_cse , mux_164_cse});
      reg_div_mgc_div_7_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_9_sg1 , else_7_else_1_if_conc_1_tmp_mut_10_sg1
          , else_7_else_1_if_conc_1_tmp_mut_11_sg1 , else_7_else_1_if_conc_1_tmp_mut_12_sg1},
          {and_994_cse , and_1000_cse , and_1007_cse , and_1015_cse , mux_164_cse});
      reg_div_mgc_div_8_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_47_sg1 ,
          mut_48_sg1 , mut_49_sg1 , mut_50_sg1}, {and_1049_cse , and_1055_cse , and_1062_cse
          , and_1070_cse , mux_171_cse});
      reg_div_mgc_div_8_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_13_sg1 , else_7_else_1_if_conc_1_tmp_mut_14_sg1
          , else_7_else_1_if_conc_1_tmp_mut_15_sg1 , else_7_else_1_if_conc_1_tmp_mut_16_sg1},
          {and_1049_cse , and_1055_cse , and_1062_cse , and_1070_cse , mux_171_cse});
      reg_div_mgc_div_9_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_51_sg1 ,
          mut_52_sg1 , mut_53_sg1 , mut_54_sg1}, {and_1104_cse , and_1110_cse , and_1117_cse
          , and_1125_cse , mux_178_cse});
      reg_div_mgc_div_9_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_17_sg1 , else_7_else_1_if_conc_1_tmp_mut_18_sg1
          , else_7_else_1_if_conc_1_tmp_mut_19_sg1 , else_7_else_1_if_conc_1_tmp_mut_20_sg1},
          {and_1104_cse , and_1110_cse , and_1117_cse , and_1125_cse , mux_178_cse});
      reg_div_mgc_div_10_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_55_sg1
          , mut_56_sg1 , mut_57_sg1 , mut_58_sg1}, {and_1159_cse , and_1165_cse ,
          and_1172_cse , and_1179_cse , mux_188_cse});
      reg_div_mgc_div_10_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_if_acc_2_itm[10:1])
          , else_7_else_1_if_conc_1_tmp_mut_21_sg1 , else_7_else_1_if_conc_1_tmp_mut_22_sg1
          , else_7_else_1_if_conc_1_tmp_mut_23_sg1 , else_7_else_1_if_conc_1_tmp_mut_24_sg1},
          {and_1159_cse , and_1165_cse , and_1172_cse , and_1179_cse , mux_188_cse});
      reg_div_mgc_div_1_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_19_sg1 ,
          mut_20_sg1 , mut_21_sg1 , mut_22_sg1}, {and_1208_cse , and_1215_cse , and_1222_cse
          , and_1230_cse , mux_198_cse});
      reg_div_mgc_div_1_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_5_sg1 , else_7_else_1_else_conc_1_tmp_mut_6_sg1
          , else_7_else_1_else_conc_1_tmp_mut_7_sg1 , else_7_else_1_else_conc_1_tmp_mut_8_sg1},
          {and_1208_cse , and_1215_cse , and_1222_cse , and_1230_cse , mux_198_cse});
      reg_div_mgc_div_2_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_23_sg1 ,
          mut_24_sg1 , mut_25_sg1 , mut_26_sg1}, {and_1264_cse , and_1270_cse , and_1277_cse
          , and_1285_cse , mux_205_cse});
      reg_div_mgc_div_2_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_9_sg1 , else_7_else_1_else_conc_1_tmp_mut_10_sg1
          , else_7_else_1_else_conc_1_tmp_mut_11_sg1 , else_7_else_1_else_conc_1_tmp_mut_12_sg1},
          {and_1264_cse , and_1270_cse , and_1277_cse , and_1285_cse , mux_205_cse});
      reg_div_mgc_div_3_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_27_sg1 ,
          mut_28_sg1 , mut_29_sg1 , mut_30_sg1}, {and_1319_cse , and_1325_cse , and_1332_cse
          , and_1340_cse , mux_212_cse});
      reg_div_mgc_div_3_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_13_sg1 , else_7_else_1_else_conc_1_tmp_mut_14_sg1
          , else_7_else_1_else_conc_1_tmp_mut_15_sg1 , else_7_else_1_else_conc_1_tmp_mut_16_sg1},
          {and_1319_cse , and_1325_cse , and_1332_cse , and_1340_cse , mux_212_cse});
      reg_div_mgc_div_4_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_31_sg1 ,
          mut_32_sg1 , mut_33_sg1 , mut_34_sg1}, {and_1374_cse , and_1380_cse , and_1387_cse
          , and_1395_cse , mux_219_cse});
      reg_div_mgc_div_4_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_17_sg1 , else_7_else_1_else_conc_1_tmp_mut_18_sg1
          , else_7_else_1_else_conc_1_tmp_mut_19_sg1 , else_7_else_1_else_conc_1_tmp_mut_20_sg1},
          {and_1374_cse , and_1380_cse , and_1387_cse , and_1395_cse , mux_219_cse});
      reg_div_mgc_div_5_b_tmp <= MUX1HOT_v_10_5_2({(acc_itm[10:1]) , mut_35_sg1 ,
          mut_36_sg1 , mut_37_sg1 , mut_38_sg1}, {and_1429_cse , and_1435_cse , and_1442_cse
          , and_1449_cse , mux_229_cse});
      reg_div_mgc_div_5_a_tmp <= MUX1HOT_v_10_5_2({(else_7_else_1_else_acc_2_itm[10:1])
          , else_7_else_1_else_conc_1_tmp_mut_21_sg1 , else_7_else_1_else_conc_1_tmp_mut_22_sg1
          , else_7_else_1_else_conc_1_tmp_mut_23_sg1 , else_7_else_1_else_conc_1_tmp_mut_24_sg1},
          {and_1429_cse , and_1435_cse , and_1442_cse , and_1449_cse , mux_229_cse});
    end
  end
  assign nl_acc_4_itm_1  = (mul_1_itm[17:8]) + conv_u2u_1_10(mul_1_itm[7]);
  assign nl_acc_5_itm_1  = conv_u2u_8_9(mul_itm[13:6]) + conv_u2u_1_9(mul_itm[5]);

  function [0:0] MUX_s_1_2_2;
    input [1:0] inputs;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[1:1];
      end
      1'b1 : begin
        result = inputs[0:0];
      end
      default : begin
        result = inputs[1:1];
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [10:0] MUX_v_11_2_2;
    input [21:0] inputs;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[21:11];
      end
      1'b1 : begin
        result = inputs[10:0];
      end
      default : begin
        result = inputs[21:11];
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function [17:0] MUX1HOT_v_18_6_2;
    input [107:0] inputs;
    input [5:0] sel;
    reg [17:0] result;
    integer i;
  begin
    result = inputs[0+:18] & {18{sel[0]}};
    for( i = 1; i < 6; i = i + 1 )
      result = result | (inputs[i*18+:18] & {18{sel[i]}});
    MUX1HOT_v_18_6_2 = result;
  end
  endfunction


  function [6:0] MUX1HOT_v_7_6_2;
    input [41:0] inputs;
    input [5:0] sel;
    reg [6:0] result;
    integer i;
  begin
    result = inputs[0+:7] & {7{sel[0]}};
    for( i = 1; i < 6; i = i + 1 )
      result = result | (inputs[i*7+:7] & {7{sel[i]}});
    MUX1HOT_v_7_6_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_6_2;
    input [35:0] inputs;
    input [5:0] sel;
    reg [5:0] result;
    integer i;
  begin
    result = inputs[0+:6] & {6{sel[0]}};
    for( i = 1; i < 6; i = i + 1 )
      result = result | (inputs[i*6+:6] & {6{sel[i]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_3_2;
    input [17:0] inputs;
    input [2:0] sel;
    reg [5:0] result;
    integer i;
  begin
    result = inputs[0+:6] & {6{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*6+:6] & {6{sel[i]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [2:0] inputs;
    input [2:0] sel;
    reg [0:0] result;
    integer i;
  begin
    result = inputs[0+:1] & {1{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*1+:1] & {1{sel[i]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [10:0] MUX1HOT_v_11_8_2;
    input [87:0] inputs;
    input [7:0] sel;
    reg [10:0] result;
    integer i;
  begin
    result = inputs[0+:11] & {11{sel[0]}};
    for( i = 1; i < 8; i = i + 1 )
      result = result | (inputs[i*11+:11] & {11{sel[i]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function [9:0] MUX1HOT_v_10_3_2;
    input [29:0] inputs;
    input [2:0] sel;
    reg [9:0] result;
    integer i;
  begin
    result = inputs[0+:10] & {10{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*10+:10] & {10{sel[i]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction


  function [17:0] MUX1HOT_v_18_3_2;
    input [53:0] inputs;
    input [2:0] sel;
    reg [17:0] result;
    integer i;
  begin
    result = inputs[0+:18] & {18{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*18+:18] & {18{sel[i]}});
    MUX1HOT_v_18_3_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [19:0] inputs;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[19:10];
      end
      1'b1 : begin
        result = inputs[9:0];
      end
      default : begin
        result = inputs[19:10];
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [13:0] inputs;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[13:7];
      end
      1'b1 : begin
        result = inputs[6:0];
      end
      default : begin
        result = inputs[13:7];
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [5:0] inputs;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[5:3];
      end
      1'b1 : begin
        result = inputs[2:0];
      end
      default : begin
        result = inputs[5:3];
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [9:0] MUX1HOT_v_10_5_2;
    input [49:0] inputs;
    input [4:0] sel;
    reg [9:0] result;
    integer i;
  begin
    result = inputs[0+:10] & {10{sel[0]}};
    for( i = 1; i < 5; i = i + 1 )
      result = result | (inputs[i*10+:10] & {10{sel[i]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function  [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function  [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function signed [2:0] conv_s2s_1_3 ;
    input signed [0:0]  vector ;
  begin
    conv_s2s_1_3 = {{2{vector[0]}}, vector};
  end
  endfunction


  function signed [2:0] conv_u2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_3 = {1'b0, vector};
  end
  endfunction


  function  [13:0] conv_u2u_10_14 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_14 = {{4{1'b0}}, vector};
  end
  endfunction


  function  [9:0] conv_u2u_1_10 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_10 = {{9{1'b0}}, vector};
  end
  endfunction


  function  [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function  [8:0] conv_u2u_1_9 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_9 = {{8{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HSVRGB
//  Generated from file(s):
//    9) $PROJECT_HOME/RGBHSV.cpp
// ------------------------------------------------------------------


module HSVRGB (
  r_rsc_z, g_rsc_z, b_rsc_z, H_OUT_rsc_z, S_OUT_rsc_z, V_OUT_rsc_z, clk, arst_n
);
  input [9:0] r_rsc_z;
  input [9:0] g_rsc_z;
  input [9:0] b_rsc_z;
  output [9:0] H_OUT_rsc_z;
  output [9:0] S_OUT_rsc_z;
  output [9:0] V_OUT_rsc_z;
  input clk;
  input arst_n;


  // Interconnect Declarations
  wire [9:0] r_rsc_mgc_in_wire_d;
  wire [9:0] g_rsc_mgc_in_wire_d;
  wire [9:0] b_rsc_mgc_in_wire_d;
  wire [9:0] H_OUT_rsc_mgc_out_stdreg_d;
  wire [9:0] S_OUT_rsc_mgc_out_stdreg_d;
  wire [9:0] V_OUT_rsc_mgc_out_stdreg_d;
  wire [29:0] div_mgc_div_a;
  wire [20:0] div_mgc_div_b;
  wire [29:0] div_mgc_div_z;
  wire [29:0] div_mgc_div_1_a;
  wire [20:0] div_mgc_div_1_b;
  wire [29:0] div_mgc_div_1_z;
  wire [29:0] div_mgc_div_2_a;
  wire [20:0] div_mgc_div_2_b;
  wire [29:0] div_mgc_div_2_z;
  wire [29:0] div_mgc_div_3_a;
  wire [20:0] div_mgc_div_3_b;
  wire [29:0] div_mgc_div_3_z;
  wire [29:0] div_mgc_div_4_a;
  wire [20:0] div_mgc_div_4_b;
  wire [29:0] div_mgc_div_4_z;
  wire [29:0] div_mgc_div_5_a;
  wire [20:0] div_mgc_div_5_b;
  wire [29:0] div_mgc_div_5_z;
  wire [29:0] div_mgc_div_6_a;
  wire [20:0] div_mgc_div_6_b;
  wire [29:0] div_mgc_div_6_z;
  wire [29:0] div_mgc_div_7_a;
  wire [20:0] div_mgc_div_7_b;
  wire [29:0] div_mgc_div_7_z;
  wire [29:0] div_mgc_div_8_a;
  wire [20:0] div_mgc_div_8_b;
  wire [29:0] div_mgc_div_8_z;
  wire [29:0] div_mgc_div_9_a;
  wire [20:0] div_mgc_div_9_b;
  wire [29:0] div_mgc_div_9_z;
  wire [29:0] div_mgc_div_10_a;
  wire [20:0] div_mgc_div_10_b;
  wire [29:0] div_mgc_div_10_z;
  wire [29:0] div_mgc_div_11_a;
  wire [20:0] div_mgc_div_11_b;
  wire [29:0] div_mgc_div_11_z;
  wire [29:0] div_mgc_div_12_a;
  wire [20:0] div_mgc_div_12_b;
  wire [29:0] div_mgc_div_12_z;
  wire [29:0] div_mgc_div_13_a;
  wire [20:0] div_mgc_div_13_b;
  wire [29:0] div_mgc_div_13_z;
  wire [29:0] div_mgc_div_14_a;
  wire [20:0] div_mgc_div_14_b;
  wire [29:0] div_mgc_div_14_z;
  wire [19:0] div_mgc_div_15_a;
  wire [9:0] div_mgc_div_15_b;
  wire [19:0] div_mgc_div_15_z;
  reg [19:0] div_mgc_div_15_z_oreg;
  wire [19:0] div_mgc_div_16_a;
  wire [9:0] div_mgc_div_16_b;
  wire [19:0] div_mgc_div_16_z;
  reg [19:0] div_mgc_div_16_z_oreg;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire #(.rscid(1),
  .width(10)) r_rsc_mgc_in_wire (
      .d(r_rsc_mgc_in_wire_d),
      .z(r_rsc_z)
    );
  mgc_in_wire #(.rscid(2),
  .width(10)) g_rsc_mgc_in_wire (
      .d(g_rsc_mgc_in_wire_d),
      .z(g_rsc_z)
    );
  mgc_in_wire #(.rscid(3),
  .width(10)) b_rsc_mgc_in_wire (
      .d(b_rsc_mgc_in_wire_d),
      .z(b_rsc_z)
    );
  mgc_out_stdreg #(.rscid(4),
  .width(10)) H_OUT_rsc_mgc_out_stdreg (
      .d(H_OUT_rsc_mgc_out_stdreg_d),
      .z(H_OUT_rsc_z)
    );
  mgc_out_stdreg #(.rscid(5),
  .width(10)) S_OUT_rsc_mgc_out_stdreg (
      .d(S_OUT_rsc_mgc_out_stdreg_d),
      .z(S_OUT_rsc_z)
    );
  mgc_out_stdreg #(.rscid(6),
  .width(10)) V_OUT_rsc_mgc_out_stdreg (
      .d(V_OUT_rsc_mgc_out_stdreg_d),
      .z(V_OUT_rsc_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div (
      .a(div_mgc_div_a),
      .b(div_mgc_div_b),
      .z(div_mgc_div_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_1 (
      .a(div_mgc_div_1_a),
      .b(div_mgc_div_1_b),
      .z(div_mgc_div_1_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_2 (
      .a(div_mgc_div_2_a),
      .b(div_mgc_div_2_b),
      .z(div_mgc_div_2_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_3 (
      .a(div_mgc_div_3_a),
      .b(div_mgc_div_3_b),
      .z(div_mgc_div_3_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_4 (
      .a(div_mgc_div_4_a),
      .b(div_mgc_div_4_b),
      .z(div_mgc_div_4_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_5 (
      .a(div_mgc_div_5_a),
      .b(div_mgc_div_5_b),
      .z(div_mgc_div_5_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_6 (
      .a(div_mgc_div_6_a),
      .b(div_mgc_div_6_b),
      .z(div_mgc_div_6_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_7 (
      .a(div_mgc_div_7_a),
      .b(div_mgc_div_7_b),
      .z(div_mgc_div_7_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_8 (
      .a(div_mgc_div_8_a),
      .b(div_mgc_div_8_b),
      .z(div_mgc_div_8_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_9 (
      .a(div_mgc_div_9_a),
      .b(div_mgc_div_9_b),
      .z(div_mgc_div_9_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_10 (
      .a(div_mgc_div_10_a),
      .b(div_mgc_div_10_b),
      .z(div_mgc_div_10_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_11 (
      .a(div_mgc_div_11_a),
      .b(div_mgc_div_11_b),
      .z(div_mgc_div_11_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_12 (
      .a(div_mgc_div_12_a),
      .b(div_mgc_div_12_b),
      .z(div_mgc_div_12_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_13 (
      .a(div_mgc_div_13_a),
      .b(div_mgc_div_13_b),
      .z(div_mgc_div_13_z)
    );
  mgc_div #(.width_a(30),
  .width_b(21),
  .signd(1)) div_mgc_div_14 (
      .a(div_mgc_div_14_a),
      .b(div_mgc_div_14_b),
      .z(div_mgc_div_14_z)
    );
  mgc_div #(.width_a(20),
  .width_b(10),
  .signd(0)) div_mgc_div_15 (
      .a(div_mgc_div_15_a),
      .b(div_mgc_div_15_b),
      .z(div_mgc_div_15_z)
    );
  mgc_div #(.width_a(20),
  .width_b(10),
  .signd(0)) div_mgc_div_16 (
      .a(div_mgc_div_16_a),
      .b(div_mgc_div_16_b),
      .z(div_mgc_div_16_z)
    );
  HSVRGB_core HSVRGB_core_inst (
      .clk(clk),
      .arst_n(arst_n),
      .r_rsc_mgc_in_wire_d(r_rsc_mgc_in_wire_d),
      .g_rsc_mgc_in_wire_d(g_rsc_mgc_in_wire_d),
      .b_rsc_mgc_in_wire_d(b_rsc_mgc_in_wire_d),
      .H_OUT_rsc_mgc_out_stdreg_d(H_OUT_rsc_mgc_out_stdreg_d),
      .S_OUT_rsc_mgc_out_stdreg_d(S_OUT_rsc_mgc_out_stdreg_d),
      .V_OUT_rsc_mgc_out_stdreg_d(V_OUT_rsc_mgc_out_stdreg_d),
      .div_mgc_div_a(div_mgc_div_a),
      .div_mgc_div_b(div_mgc_div_b),
      .div_mgc_div_z(div_mgc_div_z),
      .div_mgc_div_1_a(div_mgc_div_1_a),
      .div_mgc_div_1_b(div_mgc_div_1_b),
      .div_mgc_div_1_z(div_mgc_div_1_z),
      .div_mgc_div_2_a(div_mgc_div_2_a),
      .div_mgc_div_2_b(div_mgc_div_2_b),
      .div_mgc_div_2_z(div_mgc_div_2_z),
      .div_mgc_div_3_a(div_mgc_div_3_a),
      .div_mgc_div_3_b(div_mgc_div_3_b),
      .div_mgc_div_3_z(div_mgc_div_3_z),
      .div_mgc_div_4_a(div_mgc_div_4_a),
      .div_mgc_div_4_b(div_mgc_div_4_b),
      .div_mgc_div_4_z(div_mgc_div_4_z),
      .div_mgc_div_5_a(div_mgc_div_5_a),
      .div_mgc_div_5_b(div_mgc_div_5_b),
      .div_mgc_div_5_z(div_mgc_div_5_z),
      .div_mgc_div_6_a(div_mgc_div_6_a),
      .div_mgc_div_6_b(div_mgc_div_6_b),
      .div_mgc_div_6_z(div_mgc_div_6_z),
      .div_mgc_div_7_a(div_mgc_div_7_a),
      .div_mgc_div_7_b(div_mgc_div_7_b),
      .div_mgc_div_7_z(div_mgc_div_7_z),
      .div_mgc_div_8_a(div_mgc_div_8_a),
      .div_mgc_div_8_b(div_mgc_div_8_b),
      .div_mgc_div_8_z(div_mgc_div_8_z),
      .div_mgc_div_9_a(div_mgc_div_9_a),
      .div_mgc_div_9_b(div_mgc_div_9_b),
      .div_mgc_div_9_z(div_mgc_div_9_z),
      .div_mgc_div_10_a(div_mgc_div_10_a),
      .div_mgc_div_10_b(div_mgc_div_10_b),
      .div_mgc_div_10_z(div_mgc_div_10_z),
      .div_mgc_div_11_a(div_mgc_div_11_a),
      .div_mgc_div_11_b(div_mgc_div_11_b),
      .div_mgc_div_11_z(div_mgc_div_11_z),
      .div_mgc_div_12_a(div_mgc_div_12_a),
      .div_mgc_div_12_b(div_mgc_div_12_b),
      .div_mgc_div_12_z(div_mgc_div_12_z),
      .div_mgc_div_13_a(div_mgc_div_13_a),
      .div_mgc_div_13_b(div_mgc_div_13_b),
      .div_mgc_div_13_z(div_mgc_div_13_z),
      .div_mgc_div_14_a(div_mgc_div_14_a),
      .div_mgc_div_14_b(div_mgc_div_14_b),
      .div_mgc_div_14_z(div_mgc_div_14_z),
      .div_mgc_div_15_a(div_mgc_div_15_a),
      .div_mgc_div_15_b(div_mgc_div_15_b),
      .div_mgc_div_15_z_oreg(div_mgc_div_15_z_oreg),
      .div_mgc_div_16_a(div_mgc_div_16_a),
      .div_mgc_div_16_b(div_mgc_div_16_b),
      .div_mgc_div_16_z_oreg(div_mgc_div_16_z_oreg)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_mgc_div_15_z_oreg <= 20'b0;
      div_mgc_div_16_z_oreg <= 20'b0;
    end
    else begin
      div_mgc_div_15_z_oreg <= div_mgc_div_15_z;
      div_mgc_div_16_z_oreg <= div_mgc_div_16_z;
    end
  end
endmodule



