library verilog;
use verilog.vl_types.all;
entity TestBench_vlg_vec_tst is
end TestBench_vlg_vec_tst;
